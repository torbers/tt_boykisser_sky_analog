magic
tech sky130A
timestamp 1754386404
<< metal1 >>
rect 2996 3528 3136 3556
rect 420 3500 560 3528
rect 2912 3500 3136 3528
rect 420 3472 672 3500
rect 2856 3472 3164 3500
rect 420 3444 756 3472
rect 2772 3444 3164 3472
rect 420 3416 812 3444
rect 2716 3416 2996 3444
rect 3080 3416 3164 3444
rect 392 3332 504 3416
rect 616 3388 840 3416
rect 2660 3388 2912 3416
rect 672 3360 868 3388
rect 2604 3360 2856 3388
rect 3080 3360 3192 3416
rect 728 3332 896 3360
rect 2576 3332 2800 3360
rect 3108 3332 3192 3360
rect 392 3304 476 3332
rect 756 3304 924 3332
rect 1372 3304 1456 3332
rect 2520 3304 2744 3332
rect 364 3248 476 3304
rect 784 3276 980 3304
rect 1372 3276 1680 3304
rect 2492 3276 2688 3304
rect 3108 3276 3220 3332
rect 840 3248 1008 3276
rect 1372 3248 1764 3276
rect 2464 3248 2632 3276
rect 3136 3248 3220 3276
rect 364 3164 448 3248
rect 868 3220 1064 3248
rect 1372 3220 1848 3248
rect 2408 3220 2604 3248
rect 896 3192 1092 3220
rect 1372 3192 1484 3220
rect 1596 3192 1932 3220
rect 2380 3192 2576 3220
rect 952 3164 1120 3192
rect 1400 3164 1484 3192
rect 1708 3164 1988 3192
rect 2380 3164 2548 3192
rect 3136 3164 3248 3248
rect 336 3108 448 3164
rect 980 3136 1148 3164
rect 1008 3108 1176 3136
rect 1400 3108 1512 3164
rect 1792 3136 2044 3164
rect 2352 3136 2520 3164
rect 3164 3136 3248 3164
rect 1848 3108 2100 3136
rect 2352 3108 2492 3136
rect 336 3024 420 3108
rect 1036 3080 1204 3108
rect 1064 3052 1204 3080
rect 1428 3052 1540 3108
rect 1904 3080 2128 3108
rect 2324 3080 2436 3108
rect 1960 3052 2156 3080
rect 2296 3052 2436 3080
rect 3164 3052 3276 3136
rect 1092 3024 1232 3052
rect 1428 3024 1568 3052
rect 2016 3024 2184 3052
rect 2296 3024 2408 3052
rect 308 2968 420 3024
rect 1120 2996 1260 3024
rect 1456 2996 1596 3024
rect 2044 2996 2240 3024
rect 2268 2996 2408 3024
rect 3192 2996 3276 3052
rect 1148 2968 1288 2996
rect 1456 2968 1624 2996
rect 2100 2968 2380 2996
rect 308 2800 392 2968
rect 1176 2940 1316 2968
rect 1484 2940 1652 2968
rect 2128 2940 2380 2968
rect 3192 2940 3304 2996
rect 1204 2912 1344 2940
rect 1512 2912 1652 2940
rect 2156 2912 2352 2940
rect 1232 2884 1372 2912
rect 1540 2884 1680 2912
rect 2184 2884 2352 2912
rect 3220 2884 3304 2940
rect 1232 2856 1400 2884
rect 1456 2856 1680 2884
rect 2212 2856 2324 2884
rect 1260 2828 1680 2856
rect 1288 2800 1624 2828
rect 2240 2800 2324 2856
rect 3220 2800 3332 2884
rect 280 2744 392 2800
rect 1344 2772 1512 2800
rect 1316 2744 1484 2772
rect 280 2632 364 2744
rect 1288 2716 1456 2744
rect 3248 2716 3332 2800
rect 252 2548 364 2632
rect 1260 2688 1428 2716
rect 1260 2660 1736 2688
rect 3248 2660 3360 2716
rect 1260 2604 1820 2660
rect 1652 2576 1820 2604
rect 3276 2632 3360 2660
rect 3276 2548 3388 2632
rect 252 2464 336 2548
rect 252 2380 364 2464
rect 3276 2436 3360 2548
rect 280 2352 364 2380
rect 3248 2352 3360 2436
rect 280 2268 392 2352
rect 3248 2296 3332 2352
rect 308 2212 420 2268
rect 3220 2240 3332 2296
rect 3192 2212 3304 2240
rect 308 2184 448 2212
rect 3164 2184 3304 2212
rect 336 2128 448 2184
rect 2212 2156 2800 2184
rect 3164 2156 3276 2184
rect 2156 2128 2800 2156
rect 3136 2128 3276 2156
rect 364 2044 476 2128
rect 756 2100 1428 2128
rect 2100 2100 2800 2128
rect 3108 2100 3248 2128
rect 756 2044 1484 2100
rect 2100 2044 2436 2100
rect 2576 2044 2716 2100
rect 3080 2072 3248 2100
rect 3052 2044 3220 2072
rect 392 1988 504 2044
rect 840 2016 980 2044
rect 812 1988 980 2016
rect 420 1932 532 1988
rect 812 1960 952 1988
rect 784 1932 924 1960
rect 420 1904 560 1932
rect 448 1876 560 1904
rect 784 1876 896 1932
rect 168 1848 252 1876
rect 448 1848 588 1876
rect 168 1820 336 1848
rect 476 1820 588 1848
rect 168 1736 700 1820
rect 756 1792 868 1876
rect 1120 1792 1512 2044
rect 196 1708 308 1736
rect 756 1708 840 1792
rect 1120 1708 1484 1792
rect 2072 1708 2436 2044
rect 2604 2016 2716 2044
rect 3024 2016 3192 2044
rect 2632 1960 2744 2016
rect 3024 1988 3164 2016
rect 2968 1960 3136 1988
rect 2660 1904 2744 1960
rect 2940 1932 3444 1960
rect 2660 1820 2772 1904
rect 2912 1876 3444 1932
rect 2912 1848 3192 1876
rect 3304 1848 3444 1876
rect 2912 1820 2996 1848
rect 3276 1820 3416 1848
rect 2688 1736 2772 1820
rect 3276 1792 3388 1820
rect 3248 1764 3388 1792
rect 3220 1736 3360 1764
rect 196 1680 336 1708
rect 224 1652 364 1680
rect 252 1624 392 1652
rect 756 1624 868 1708
rect 1148 1652 1456 1708
rect 2100 1652 2408 1708
rect 2660 1652 2772 1736
rect 3192 1708 3332 1736
rect 3164 1680 3304 1708
rect 3136 1652 3276 1680
rect 1176 1624 1428 1652
rect 2128 1624 2380 1652
rect 252 1596 420 1624
rect 280 1568 448 1596
rect 308 1540 476 1568
rect 784 1540 896 1624
rect 1176 1596 1400 1624
rect 2184 1596 2324 1624
rect 2660 1596 2744 1652
rect 3108 1624 3276 1652
rect 3080 1596 3248 1624
rect 1204 1568 1372 1596
rect 3052 1568 3220 1596
rect 336 1512 504 1540
rect 812 1512 896 1540
rect 364 1484 532 1512
rect 672 1484 784 1512
rect 1568 1484 1792 1568
rect 3024 1540 3192 1568
rect 2548 1512 2660 1540
rect 2492 1484 2660 1512
rect 2744 1484 2856 1512
rect 392 1456 532 1484
rect 644 1456 812 1484
rect 2464 1456 2660 1484
rect 2716 1456 2856 1484
rect 3024 1484 3164 1540
rect 3024 1456 3192 1484
rect 420 1428 532 1456
rect 588 1428 812 1456
rect 924 1428 1008 1456
rect 2436 1428 2856 1456
rect 3052 1428 3220 1456
rect 392 1400 532 1428
rect 560 1400 840 1428
rect 896 1400 1008 1428
rect 392 1372 504 1400
rect 364 1344 504 1372
rect 560 1372 700 1400
rect 560 1344 672 1372
rect 728 1344 1008 1400
rect 2408 1400 2828 1428
rect 3080 1400 3248 1428
rect 2408 1372 2548 1400
rect 2576 1372 2800 1400
rect 3108 1372 3248 1400
rect 2072 1344 2156 1372
rect 2408 1344 2520 1372
rect 2576 1344 2744 1372
rect 3136 1344 3276 1372
rect 364 1316 476 1344
rect 336 1288 476 1316
rect 756 1316 980 1344
rect 1708 1316 1792 1344
rect 2016 1316 2156 1344
rect 756 1288 924 1316
rect 1680 1288 1820 1316
rect 1988 1288 2156 1316
rect 2576 1316 2716 1344
rect 2576 1288 2688 1316
rect 3164 1288 3304 1344
rect 336 1232 448 1288
rect 1652 1260 2156 1288
rect 1400 1232 1540 1260
rect 1596 1232 2100 1260
rect 3192 1232 3332 1288
rect 336 1148 420 1232
rect 1400 1204 2072 1232
rect 3136 1204 3332 1232
rect 1400 1176 1736 1204
rect 1820 1176 1988 1204
rect 2688 1176 2800 1204
rect 3080 1176 3304 1204
rect 1456 1148 1680 1176
rect 2660 1148 2800 1176
rect 2912 1148 3276 1176
rect 336 1120 504 1148
rect 644 1120 868 1148
rect 2632 1120 3220 1148
rect 336 1092 924 1120
rect 2576 1092 2772 1120
rect 2800 1092 3136 1120
rect 336 1064 952 1092
rect 2520 1064 2744 1092
rect 2800 1064 2996 1092
rect 420 1036 728 1064
rect 784 1036 1008 1064
rect 2464 1036 2716 1064
rect 840 1008 1064 1036
rect 2380 1008 2660 1036
rect 868 980 1288 1008
rect 2296 980 2604 1008
rect 924 952 1344 980
rect 2296 952 2520 980
rect 980 924 1512 952
rect 2296 924 2436 952
rect 1036 896 1148 924
rect 1204 896 1512 924
rect 1036 868 1176 896
rect 1288 868 1512 896
rect 1064 840 1176 868
rect 2408 840 2520 896
rect 1064 812 1204 840
rect 2408 812 2548 840
rect 1092 784 1232 812
rect 1092 756 1260 784
rect 2436 756 2576 812
rect 1120 728 1288 756
rect 2464 728 2576 756
rect 1148 700 1316 728
rect 1176 672 1316 700
rect 2492 672 2604 728
rect 1204 644 1316 672
rect 1176 588 1316 644
rect 2520 588 2632 672
rect 1148 560 1288 588
rect 2548 560 2632 588
rect 1120 532 1260 560
rect 1092 504 1232 532
rect 1064 476 1232 504
rect 2548 476 2660 560
rect 1064 448 1372 476
rect 1064 392 1400 448
rect 2576 392 2688 476
rect 1260 364 1400 392
rect 2604 364 2688 392
rect 1260 308 1372 364
rect 2604 308 2716 364
rect 1232 252 1344 308
rect 2632 252 2716 308
rect 1232 224 1316 252
rect 1204 168 1316 224
rect 2632 168 2744 252
rect 1204 28 1288 168
rect 2660 28 2744 168
<< obsm1 >>
rect 0 3556 3584 3584
rect 0 3528 2996 3556
rect 0 3416 420 3528
rect 560 3500 2912 3528
rect 3136 3500 3584 3556
rect 672 3472 2856 3500
rect 756 3444 2772 3472
rect 812 3416 2716 3444
rect 2996 3416 3080 3444
rect 3164 3416 3584 3500
rect 0 3304 392 3416
rect 504 3388 616 3416
rect 840 3388 2660 3416
rect 2912 3388 3080 3416
rect 504 3360 672 3388
rect 868 3360 2604 3388
rect 2856 3360 3080 3388
rect 504 3332 728 3360
rect 896 3332 2576 3360
rect 2800 3332 3108 3360
rect 3192 3332 3584 3416
rect 476 3304 756 3332
rect 924 3304 1372 3332
rect 1456 3304 2520 3332
rect 2744 3304 3108 3332
rect 0 3164 364 3304
rect 476 3276 784 3304
rect 980 3276 1372 3304
rect 1680 3276 2492 3304
rect 2688 3276 3108 3304
rect 476 3248 840 3276
rect 1008 3248 1372 3276
rect 1764 3248 2464 3276
rect 2632 3248 3136 3276
rect 3220 3248 3584 3332
rect 448 3220 868 3248
rect 1064 3220 1372 3248
rect 1848 3220 2408 3248
rect 2604 3220 3136 3248
rect 448 3192 896 3220
rect 1092 3192 1372 3220
rect 1484 3192 1596 3220
rect 1932 3192 2380 3220
rect 2576 3192 3136 3220
rect 448 3164 952 3192
rect 1120 3164 1400 3192
rect 1484 3164 1708 3192
rect 1988 3164 2380 3192
rect 2548 3164 3136 3192
rect 0 3024 336 3164
rect 448 3136 980 3164
rect 1148 3136 1400 3164
rect 448 3108 1008 3136
rect 1176 3108 1400 3136
rect 1512 3136 1792 3164
rect 2044 3136 2352 3164
rect 2520 3136 3164 3164
rect 3248 3136 3584 3248
rect 1512 3108 1848 3136
rect 2100 3108 2352 3136
rect 2492 3108 3164 3136
rect 420 3080 1036 3108
rect 420 3052 1064 3080
rect 1204 3052 1428 3108
rect 1540 3080 1904 3108
rect 2128 3080 2324 3108
rect 1540 3052 1960 3080
rect 2156 3052 2296 3080
rect 2436 3052 3164 3108
rect 420 3024 1092 3052
rect 1232 3024 1428 3052
rect 1568 3024 2016 3052
rect 2184 3024 2296 3052
rect 0 2800 308 3024
rect 420 2996 1120 3024
rect 1260 2996 1456 3024
rect 1596 2996 2044 3024
rect 2240 2996 2268 3024
rect 2408 2996 3192 3052
rect 3276 2996 3584 3136
rect 420 2968 1148 2996
rect 1288 2968 1456 2996
rect 1624 2968 2100 2996
rect 392 2940 1176 2968
rect 1316 2940 1484 2968
rect 1652 2940 2128 2968
rect 2380 2940 3192 2996
rect 392 2912 1204 2940
rect 1344 2912 1512 2940
rect 1652 2912 2156 2940
rect 392 2856 1232 2912
rect 1372 2884 1540 2912
rect 1680 2884 2184 2912
rect 2352 2884 3220 2940
rect 3304 2884 3584 2996
rect 1400 2856 1456 2884
rect 1680 2856 2212 2884
rect 392 2828 1260 2856
rect 1680 2828 2240 2856
rect 392 2800 1288 2828
rect 1624 2800 2240 2828
rect 2324 2800 3220 2884
rect 0 2632 280 2800
rect 392 2772 1344 2800
rect 1512 2772 3248 2800
rect 392 2744 1316 2772
rect 1484 2744 3248 2772
rect 364 2716 1288 2744
rect 1456 2716 3248 2744
rect 3332 2716 3584 2884
rect 0 2380 252 2632
rect 364 2604 1260 2716
rect 1428 2688 3248 2716
rect 1736 2660 3248 2688
rect 364 2576 1652 2604
rect 1820 2576 3276 2660
rect 3360 2632 3584 2716
rect 364 2548 3276 2576
rect 3388 2548 3584 2632
rect 336 2464 3276 2548
rect 364 2436 3276 2464
rect 0 2268 280 2380
rect 364 2352 3248 2436
rect 3360 2352 3584 2548
rect 392 2296 3248 2352
rect 392 2268 3220 2296
rect 0 2184 308 2268
rect 420 2240 3220 2268
rect 3332 2240 3584 2352
rect 420 2212 3192 2240
rect 448 2184 3164 2212
rect 3304 2184 3584 2240
rect 0 2128 336 2184
rect 448 2156 2212 2184
rect 2800 2156 3164 2184
rect 448 2128 2156 2156
rect 2800 2128 3136 2156
rect 3276 2128 3584 2184
rect 0 2044 364 2128
rect 476 2044 756 2128
rect 1428 2100 2100 2128
rect 2800 2100 3108 2128
rect 1484 2044 2100 2100
rect 2436 2044 2576 2100
rect 2716 2072 3080 2100
rect 3248 2072 3584 2128
rect 2716 2044 3052 2072
rect 3220 2044 3584 2072
rect 0 1988 392 2044
rect 504 2016 840 2044
rect 504 1988 812 2016
rect 980 1988 1120 2044
rect 0 1904 420 1988
rect 532 1960 812 1988
rect 952 1960 1120 1988
rect 532 1932 784 1960
rect 924 1932 1120 1960
rect 0 1876 448 1904
rect 560 1876 784 1932
rect 896 1876 1120 1932
rect 0 1736 168 1876
rect 252 1848 448 1876
rect 336 1820 476 1848
rect 588 1820 756 1876
rect 700 1736 756 1820
rect 868 1792 1120 1876
rect 1512 1792 2072 2044
rect 0 1680 196 1736
rect 308 1708 756 1736
rect 840 1708 1120 1792
rect 1484 1708 2072 1792
rect 2436 2016 2604 2044
rect 2716 2016 3024 2044
rect 3192 2016 3584 2044
rect 2436 1960 2632 2016
rect 2744 1988 3024 2016
rect 3164 1988 3584 2016
rect 2744 1960 2968 1988
rect 3136 1960 3584 1988
rect 2436 1820 2660 1960
rect 2744 1932 2940 1960
rect 2744 1904 2912 1932
rect 2772 1820 2912 1904
rect 3192 1848 3304 1876
rect 3444 1848 3584 1960
rect 2996 1820 3276 1848
rect 3416 1820 3584 1848
rect 2436 1736 2688 1820
rect 2772 1792 3276 1820
rect 2772 1764 3248 1792
rect 3388 1764 3584 1820
rect 2772 1736 3220 1764
rect 3360 1736 3584 1764
rect 2436 1708 2660 1736
rect 336 1680 756 1708
rect 0 1652 224 1680
rect 364 1652 756 1680
rect 0 1596 252 1652
rect 392 1624 756 1652
rect 868 1652 1148 1708
rect 1456 1652 2100 1708
rect 2408 1652 2660 1708
rect 2772 1708 3192 1736
rect 3332 1708 3584 1736
rect 2772 1680 3164 1708
rect 3304 1680 3584 1708
rect 2772 1652 3136 1680
rect 868 1624 1176 1652
rect 1428 1624 2128 1652
rect 2380 1624 2660 1652
rect 420 1596 784 1624
rect 0 1568 280 1596
rect 448 1568 784 1596
rect 0 1540 308 1568
rect 476 1540 784 1568
rect 896 1596 1176 1624
rect 1400 1596 2184 1624
rect 2324 1596 2660 1624
rect 2744 1624 3108 1652
rect 3276 1624 3584 1680
rect 2744 1596 3080 1624
rect 3248 1596 3584 1624
rect 896 1568 1204 1596
rect 1372 1568 3052 1596
rect 3220 1568 3584 1596
rect 0 1512 336 1540
rect 504 1512 812 1540
rect 896 1512 1568 1568
rect 0 1484 364 1512
rect 532 1484 672 1512
rect 784 1484 1568 1512
rect 1792 1540 3024 1568
rect 3192 1540 3584 1568
rect 1792 1512 2548 1540
rect 2660 1512 3024 1540
rect 1792 1484 2492 1512
rect 2660 1484 2744 1512
rect 0 1456 392 1484
rect 532 1456 644 1484
rect 812 1456 2464 1484
rect 2660 1456 2716 1484
rect 2856 1456 3024 1512
rect 3164 1484 3584 1540
rect 3192 1456 3584 1484
rect 0 1428 420 1456
rect 532 1428 588 1456
rect 812 1428 924 1456
rect 1008 1428 2436 1456
rect 2856 1428 3052 1456
rect 3220 1428 3584 1456
rect 0 1372 392 1428
rect 532 1400 560 1428
rect 840 1400 896 1428
rect 0 1316 364 1372
rect 504 1344 560 1400
rect 700 1372 728 1400
rect 672 1344 728 1372
rect 1008 1372 2408 1428
rect 2828 1400 3080 1428
rect 2548 1372 2576 1400
rect 2800 1372 3108 1400
rect 3248 1372 3584 1428
rect 1008 1344 2072 1372
rect 2156 1344 2408 1372
rect 2520 1344 2576 1372
rect 2744 1344 3136 1372
rect 3276 1344 3584 1372
rect 0 1064 336 1316
rect 476 1288 756 1344
rect 980 1316 1708 1344
rect 1792 1316 2016 1344
rect 924 1288 1680 1316
rect 1820 1288 1988 1316
rect 2156 1288 2576 1344
rect 2716 1316 3164 1344
rect 2688 1288 3164 1316
rect 3304 1288 3584 1344
rect 448 1260 1652 1288
rect 2156 1260 3192 1288
rect 448 1232 1400 1260
rect 1540 1232 1596 1260
rect 2100 1232 3192 1260
rect 420 1176 1400 1232
rect 2072 1204 3136 1232
rect 3332 1204 3584 1288
rect 1736 1176 1820 1204
rect 1988 1176 2688 1204
rect 2800 1176 3080 1204
rect 3304 1176 3584 1204
rect 420 1148 1456 1176
rect 1680 1148 2660 1176
rect 2800 1148 2912 1176
rect 3276 1148 3584 1176
rect 504 1120 644 1148
rect 868 1120 2632 1148
rect 3220 1120 3584 1148
rect 924 1092 2576 1120
rect 2772 1092 2800 1120
rect 3136 1092 3584 1120
rect 952 1064 2520 1092
rect 2744 1064 2800 1092
rect 2996 1064 3584 1092
rect 0 1036 420 1064
rect 728 1036 784 1064
rect 1008 1036 2464 1064
rect 2716 1036 3584 1064
rect 0 1008 840 1036
rect 1064 1008 2380 1036
rect 2660 1008 3584 1036
rect 0 980 868 1008
rect 1288 980 2296 1008
rect 2604 980 3584 1008
rect 0 952 924 980
rect 1344 952 2296 980
rect 2520 952 3584 980
rect 0 924 980 952
rect 1512 924 2296 952
rect 2436 924 3584 952
rect 0 868 1036 924
rect 1148 896 1204 924
rect 1512 896 3584 924
rect 1176 868 1288 896
rect 1512 868 2408 896
rect 0 812 1064 868
rect 1176 840 2408 868
rect 2520 840 3584 896
rect 1204 812 2408 840
rect 2548 812 3584 840
rect 0 756 1092 812
rect 1232 784 2436 812
rect 1260 756 2436 784
rect 0 728 1120 756
rect 1288 728 2464 756
rect 2576 728 3584 812
rect 0 700 1148 728
rect 0 672 1176 700
rect 1316 672 2492 728
rect 2604 672 3584 728
rect 0 644 1204 672
rect 0 588 1176 644
rect 1316 588 2520 672
rect 0 560 1148 588
rect 1288 560 2548 588
rect 2632 560 3584 672
rect 0 532 1120 560
rect 1260 532 2548 560
rect 0 504 1092 532
rect 0 392 1064 504
rect 1232 476 2548 532
rect 2660 476 3584 560
rect 1372 448 2576 476
rect 1400 392 2576 448
rect 0 308 1260 392
rect 1400 364 2604 392
rect 2688 364 3584 476
rect 1372 308 2604 364
rect 0 224 1232 308
rect 1344 252 2632 308
rect 2716 252 3584 364
rect 0 28 1204 224
rect 1316 168 2632 252
rect 1288 28 2660 168
rect 2744 28 3584 252
rect 0 0 3584 28
<< metal2 >>
rect 2996 3528 3136 3556
rect 420 3500 560 3528
rect 2912 3500 3136 3528
rect 420 3472 672 3500
rect 2856 3472 3164 3500
rect 420 3444 756 3472
rect 2772 3444 3164 3472
rect 420 3416 812 3444
rect 2716 3416 2996 3444
rect 3080 3416 3164 3444
rect 392 3332 504 3416
rect 616 3388 840 3416
rect 2660 3388 2912 3416
rect 672 3360 868 3388
rect 2604 3360 2856 3388
rect 3080 3360 3192 3416
rect 728 3332 896 3360
rect 2576 3332 2800 3360
rect 3108 3332 3192 3360
rect 392 3304 476 3332
rect 756 3304 924 3332
rect 1372 3304 1456 3332
rect 2520 3304 2744 3332
rect 364 3248 476 3304
rect 784 3276 980 3304
rect 1372 3276 1680 3304
rect 2492 3276 2688 3304
rect 3108 3276 3220 3332
rect 840 3248 1008 3276
rect 1372 3248 1764 3276
rect 2464 3248 2632 3276
rect 3136 3248 3220 3276
rect 364 3164 448 3248
rect 868 3220 1064 3248
rect 1372 3220 1848 3248
rect 2408 3220 2604 3248
rect 896 3192 1092 3220
rect 1372 3192 1484 3220
rect 1596 3192 1932 3220
rect 2380 3192 2576 3220
rect 952 3164 1120 3192
rect 1400 3164 1484 3192
rect 1708 3164 1988 3192
rect 2380 3164 2548 3192
rect 3136 3164 3248 3248
rect 336 3108 448 3164
rect 980 3136 1148 3164
rect 1008 3108 1176 3136
rect 1400 3108 1512 3164
rect 1792 3136 2044 3164
rect 2352 3136 2520 3164
rect 3164 3136 3248 3164
rect 1848 3108 2100 3136
rect 2352 3108 2492 3136
rect 336 3024 420 3108
rect 1036 3080 1204 3108
rect 1064 3052 1204 3080
rect 1428 3052 1540 3108
rect 1904 3080 2128 3108
rect 2324 3080 2436 3108
rect 1960 3052 2156 3080
rect 2296 3052 2436 3080
rect 3164 3052 3276 3136
rect 1092 3024 1232 3052
rect 1428 3024 1568 3052
rect 2016 3024 2184 3052
rect 2296 3024 2408 3052
rect 308 2968 420 3024
rect 1120 2996 1260 3024
rect 1456 2996 1596 3024
rect 2044 2996 2240 3024
rect 2268 2996 2408 3024
rect 3192 2996 3276 3052
rect 1148 2968 1288 2996
rect 1456 2968 1624 2996
rect 2100 2968 2380 2996
rect 308 2800 392 2968
rect 1176 2940 1316 2968
rect 1484 2940 1652 2968
rect 2128 2940 2380 2968
rect 3192 2940 3304 2996
rect 1204 2912 1344 2940
rect 1512 2912 1652 2940
rect 2156 2912 2352 2940
rect 1232 2884 1372 2912
rect 1540 2884 1680 2912
rect 2184 2884 2352 2912
rect 3220 2884 3304 2940
rect 1232 2856 1400 2884
rect 1456 2856 1680 2884
rect 2212 2856 2324 2884
rect 1260 2828 1680 2856
rect 1288 2800 1624 2828
rect 2240 2800 2324 2856
rect 3220 2800 3332 2884
rect 280 2744 392 2800
rect 1344 2772 1512 2800
rect 1316 2744 1484 2772
rect 280 2632 364 2744
rect 1288 2716 1456 2744
rect 3248 2716 3332 2800
rect 252 2548 364 2632
rect 1260 2688 1428 2716
rect 1260 2660 1736 2688
rect 3248 2660 3360 2716
rect 1260 2604 1820 2660
rect 1652 2576 1820 2604
rect 3276 2632 3360 2660
rect 3276 2548 3388 2632
rect 252 2464 336 2548
rect 252 2380 364 2464
rect 3276 2436 3360 2548
rect 280 2352 364 2380
rect 3248 2352 3360 2436
rect 280 2268 392 2352
rect 3248 2296 3332 2352
rect 308 2212 420 2268
rect 3220 2240 3332 2296
rect 3192 2212 3304 2240
rect 308 2184 448 2212
rect 3164 2184 3304 2212
rect 336 2128 448 2184
rect 2212 2156 2800 2184
rect 3164 2156 3276 2184
rect 2156 2128 2800 2156
rect 3136 2128 3276 2156
rect 364 2044 476 2128
rect 756 2100 1428 2128
rect 2100 2100 2800 2128
rect 3108 2100 3248 2128
rect 756 2044 1484 2100
rect 2100 2044 2436 2100
rect 2576 2044 2716 2100
rect 3080 2072 3248 2100
rect 3052 2044 3220 2072
rect 392 1988 504 2044
rect 840 2016 980 2044
rect 812 1988 980 2016
rect 420 1932 532 1988
rect 812 1960 952 1988
rect 784 1932 924 1960
rect 420 1904 560 1932
rect 448 1876 560 1904
rect 784 1876 896 1932
rect 168 1848 252 1876
rect 448 1848 588 1876
rect 168 1820 336 1848
rect 476 1820 588 1848
rect 168 1736 700 1820
rect 756 1792 868 1876
rect 1120 1792 1512 2044
rect 196 1708 308 1736
rect 756 1708 840 1792
rect 1120 1708 1484 1792
rect 2072 1708 2436 2044
rect 2604 2016 2716 2044
rect 3024 2016 3192 2044
rect 2632 1960 2744 2016
rect 3024 1988 3164 2016
rect 2968 1960 3136 1988
rect 2660 1904 2744 1960
rect 2940 1932 3444 1960
rect 2660 1820 2772 1904
rect 2912 1876 3444 1932
rect 2912 1848 3192 1876
rect 3304 1848 3444 1876
rect 2912 1820 2996 1848
rect 3276 1820 3416 1848
rect 2688 1736 2772 1820
rect 3276 1792 3388 1820
rect 3248 1764 3388 1792
rect 3220 1736 3360 1764
rect 196 1680 336 1708
rect 224 1652 364 1680
rect 252 1624 392 1652
rect 756 1624 868 1708
rect 1148 1652 1456 1708
rect 2100 1652 2408 1708
rect 2660 1652 2772 1736
rect 3192 1708 3332 1736
rect 3164 1680 3304 1708
rect 3136 1652 3276 1680
rect 1176 1624 1428 1652
rect 2128 1624 2380 1652
rect 252 1596 420 1624
rect 280 1568 448 1596
rect 308 1540 476 1568
rect 784 1540 896 1624
rect 1176 1596 1400 1624
rect 2184 1596 2324 1624
rect 2660 1596 2744 1652
rect 3108 1624 3276 1652
rect 3080 1596 3248 1624
rect 1204 1568 1372 1596
rect 3052 1568 3220 1596
rect 336 1512 504 1540
rect 812 1512 896 1540
rect 364 1484 532 1512
rect 672 1484 784 1512
rect 1568 1484 1792 1568
rect 3024 1540 3192 1568
rect 2548 1512 2660 1540
rect 2492 1484 2660 1512
rect 2744 1484 2856 1512
rect 392 1456 532 1484
rect 644 1456 812 1484
rect 2464 1456 2660 1484
rect 2716 1456 2856 1484
rect 3024 1484 3164 1540
rect 3024 1456 3192 1484
rect 420 1428 532 1456
rect 588 1428 812 1456
rect 924 1428 1008 1456
rect 2436 1428 2856 1456
rect 3052 1428 3220 1456
rect 392 1400 532 1428
rect 560 1400 840 1428
rect 896 1400 1008 1428
rect 392 1372 504 1400
rect 364 1344 504 1372
rect 560 1372 700 1400
rect 560 1344 672 1372
rect 728 1344 1008 1400
rect 2408 1400 2828 1428
rect 3080 1400 3248 1428
rect 2408 1372 2548 1400
rect 2576 1372 2800 1400
rect 3108 1372 3248 1400
rect 2072 1344 2156 1372
rect 2408 1344 2520 1372
rect 2576 1344 2744 1372
rect 3136 1344 3276 1372
rect 364 1316 476 1344
rect 336 1288 476 1316
rect 756 1316 980 1344
rect 1708 1316 1792 1344
rect 2016 1316 2156 1344
rect 756 1288 924 1316
rect 1680 1288 1820 1316
rect 1988 1288 2156 1316
rect 2576 1316 2716 1344
rect 2576 1288 2688 1316
rect 3164 1288 3304 1344
rect 336 1232 448 1288
rect 1652 1260 2156 1288
rect 1400 1232 1540 1260
rect 1596 1232 2100 1260
rect 3192 1232 3332 1288
rect 336 1148 420 1232
rect 1400 1204 2072 1232
rect 3136 1204 3332 1232
rect 1400 1176 1736 1204
rect 1820 1176 1988 1204
rect 2688 1176 2800 1204
rect 3080 1176 3304 1204
rect 1456 1148 1680 1176
rect 2660 1148 2800 1176
rect 2912 1148 3276 1176
rect 336 1120 504 1148
rect 644 1120 868 1148
rect 2632 1120 3220 1148
rect 336 1092 924 1120
rect 2576 1092 2772 1120
rect 2800 1092 3136 1120
rect 336 1064 952 1092
rect 2520 1064 2744 1092
rect 2800 1064 2996 1092
rect 420 1036 728 1064
rect 784 1036 1008 1064
rect 2464 1036 2716 1064
rect 840 1008 1064 1036
rect 2380 1008 2660 1036
rect 868 980 1288 1008
rect 2296 980 2604 1008
rect 924 952 1344 980
rect 2296 952 2520 980
rect 980 924 1512 952
rect 2296 924 2436 952
rect 1036 896 1148 924
rect 1204 896 1512 924
rect 1036 868 1176 896
rect 1288 868 1512 896
rect 1064 840 1176 868
rect 2408 840 2520 896
rect 1064 812 1204 840
rect 2408 812 2548 840
rect 1092 784 1232 812
rect 1092 756 1260 784
rect 2436 756 2576 812
rect 1120 728 1288 756
rect 2464 728 2576 756
rect 1148 700 1316 728
rect 1176 672 1316 700
rect 2492 672 2604 728
rect 1204 644 1316 672
rect 1176 588 1316 644
rect 2520 588 2632 672
rect 1148 560 1288 588
rect 2548 560 2632 588
rect 1120 532 1260 560
rect 1092 504 1232 532
rect 1064 476 1232 504
rect 2548 476 2660 560
rect 1064 448 1372 476
rect 1064 392 1400 448
rect 2576 392 2688 476
rect 1260 364 1400 392
rect 2604 364 2688 392
rect 1260 308 1372 364
rect 2604 308 2716 364
rect 1232 252 1344 308
rect 2632 252 2716 308
rect 1232 224 1316 252
rect 1204 168 1316 224
rect 2632 168 2744 252
rect 1204 28 1288 168
rect 2660 28 2744 168
<< obsm2 >>
rect 0 3556 3584 3584
rect 0 3528 2996 3556
rect 0 3416 420 3528
rect 560 3500 2912 3528
rect 3136 3500 3584 3556
rect 672 3472 2856 3500
rect 756 3444 2772 3472
rect 812 3416 2716 3444
rect 2996 3416 3080 3444
rect 3164 3416 3584 3500
rect 0 3304 392 3416
rect 504 3388 616 3416
rect 840 3388 2660 3416
rect 2912 3388 3080 3416
rect 504 3360 672 3388
rect 868 3360 2604 3388
rect 2856 3360 3080 3388
rect 504 3332 728 3360
rect 896 3332 2576 3360
rect 2800 3332 3108 3360
rect 3192 3332 3584 3416
rect 476 3304 756 3332
rect 924 3304 1372 3332
rect 1456 3304 2520 3332
rect 2744 3304 3108 3332
rect 0 3164 364 3304
rect 476 3276 784 3304
rect 980 3276 1372 3304
rect 1680 3276 2492 3304
rect 2688 3276 3108 3304
rect 476 3248 840 3276
rect 1008 3248 1372 3276
rect 1764 3248 2464 3276
rect 2632 3248 3136 3276
rect 3220 3248 3584 3332
rect 448 3220 868 3248
rect 1064 3220 1372 3248
rect 1848 3220 2408 3248
rect 2604 3220 3136 3248
rect 448 3192 896 3220
rect 1092 3192 1372 3220
rect 1484 3192 1596 3220
rect 1932 3192 2380 3220
rect 2576 3192 3136 3220
rect 448 3164 952 3192
rect 1120 3164 1400 3192
rect 1484 3164 1708 3192
rect 1988 3164 2380 3192
rect 2548 3164 3136 3192
rect 0 3024 336 3164
rect 448 3136 980 3164
rect 1148 3136 1400 3164
rect 448 3108 1008 3136
rect 1176 3108 1400 3136
rect 1512 3136 1792 3164
rect 2044 3136 2352 3164
rect 2520 3136 3164 3164
rect 3248 3136 3584 3248
rect 1512 3108 1848 3136
rect 2100 3108 2352 3136
rect 2492 3108 3164 3136
rect 420 3080 1036 3108
rect 420 3052 1064 3080
rect 1204 3052 1428 3108
rect 1540 3080 1904 3108
rect 2128 3080 2324 3108
rect 1540 3052 1960 3080
rect 2156 3052 2296 3080
rect 2436 3052 3164 3108
rect 420 3024 1092 3052
rect 1232 3024 1428 3052
rect 1568 3024 2016 3052
rect 2184 3024 2296 3052
rect 0 2800 308 3024
rect 420 2996 1120 3024
rect 1260 2996 1456 3024
rect 1596 2996 2044 3024
rect 2240 2996 2268 3024
rect 2408 2996 3192 3052
rect 3276 2996 3584 3136
rect 420 2968 1148 2996
rect 1288 2968 1456 2996
rect 1624 2968 2100 2996
rect 392 2940 1176 2968
rect 1316 2940 1484 2968
rect 1652 2940 2128 2968
rect 2380 2940 3192 2996
rect 392 2912 1204 2940
rect 1344 2912 1512 2940
rect 1652 2912 2156 2940
rect 392 2856 1232 2912
rect 1372 2884 1540 2912
rect 1680 2884 2184 2912
rect 2352 2884 3220 2940
rect 3304 2884 3584 2996
rect 1400 2856 1456 2884
rect 1680 2856 2212 2884
rect 392 2828 1260 2856
rect 1680 2828 2240 2856
rect 392 2800 1288 2828
rect 1624 2800 2240 2828
rect 2324 2800 3220 2884
rect 0 2632 280 2800
rect 392 2772 1344 2800
rect 1512 2772 3248 2800
rect 392 2744 1316 2772
rect 1484 2744 3248 2772
rect 364 2716 1288 2744
rect 1456 2716 3248 2744
rect 3332 2716 3584 2884
rect 0 2380 252 2632
rect 364 2604 1260 2716
rect 1428 2688 3248 2716
rect 1736 2660 3248 2688
rect 364 2576 1652 2604
rect 1820 2576 3276 2660
rect 3360 2632 3584 2716
rect 364 2548 3276 2576
rect 3388 2548 3584 2632
rect 336 2464 3276 2548
rect 364 2436 3276 2464
rect 0 2268 280 2380
rect 364 2352 3248 2436
rect 3360 2352 3584 2548
rect 392 2296 3248 2352
rect 392 2268 3220 2296
rect 0 2184 308 2268
rect 420 2240 3220 2268
rect 3332 2240 3584 2352
rect 420 2212 3192 2240
rect 448 2184 3164 2212
rect 3304 2184 3584 2240
rect 0 2128 336 2184
rect 448 2156 2212 2184
rect 2800 2156 3164 2184
rect 448 2128 2156 2156
rect 2800 2128 3136 2156
rect 3276 2128 3584 2184
rect 0 2044 364 2128
rect 476 2044 756 2128
rect 1428 2100 2100 2128
rect 2800 2100 3108 2128
rect 1484 2044 2100 2100
rect 2436 2044 2576 2100
rect 2716 2072 3080 2100
rect 3248 2072 3584 2128
rect 2716 2044 3052 2072
rect 3220 2044 3584 2072
rect 0 1988 392 2044
rect 504 2016 840 2044
rect 504 1988 812 2016
rect 980 1988 1120 2044
rect 0 1904 420 1988
rect 532 1960 812 1988
rect 952 1960 1120 1988
rect 532 1932 784 1960
rect 924 1932 1120 1960
rect 0 1876 448 1904
rect 560 1876 784 1932
rect 896 1876 1120 1932
rect 0 1736 168 1876
rect 252 1848 448 1876
rect 336 1820 476 1848
rect 588 1820 756 1876
rect 700 1736 756 1820
rect 868 1792 1120 1876
rect 1512 1792 2072 2044
rect 0 1680 196 1736
rect 308 1708 756 1736
rect 840 1708 1120 1792
rect 1484 1708 2072 1792
rect 2436 2016 2604 2044
rect 2716 2016 3024 2044
rect 3192 2016 3584 2044
rect 2436 1960 2632 2016
rect 2744 1988 3024 2016
rect 3164 1988 3584 2016
rect 2744 1960 2968 1988
rect 3136 1960 3584 1988
rect 2436 1820 2660 1960
rect 2744 1932 2940 1960
rect 2744 1904 2912 1932
rect 2772 1820 2912 1904
rect 3192 1848 3304 1876
rect 3444 1848 3584 1960
rect 2996 1820 3276 1848
rect 3416 1820 3584 1848
rect 2436 1736 2688 1820
rect 2772 1792 3276 1820
rect 2772 1764 3248 1792
rect 3388 1764 3584 1820
rect 2772 1736 3220 1764
rect 3360 1736 3584 1764
rect 2436 1708 2660 1736
rect 336 1680 756 1708
rect 0 1652 224 1680
rect 364 1652 756 1680
rect 0 1596 252 1652
rect 392 1624 756 1652
rect 868 1652 1148 1708
rect 1456 1652 2100 1708
rect 2408 1652 2660 1708
rect 2772 1708 3192 1736
rect 3332 1708 3584 1736
rect 2772 1680 3164 1708
rect 3304 1680 3584 1708
rect 2772 1652 3136 1680
rect 868 1624 1176 1652
rect 1428 1624 2128 1652
rect 2380 1624 2660 1652
rect 420 1596 784 1624
rect 0 1568 280 1596
rect 448 1568 784 1596
rect 0 1540 308 1568
rect 476 1540 784 1568
rect 896 1596 1176 1624
rect 1400 1596 2184 1624
rect 2324 1596 2660 1624
rect 2744 1624 3108 1652
rect 3276 1624 3584 1680
rect 2744 1596 3080 1624
rect 3248 1596 3584 1624
rect 896 1568 1204 1596
rect 1372 1568 3052 1596
rect 3220 1568 3584 1596
rect 0 1512 336 1540
rect 504 1512 812 1540
rect 896 1512 1568 1568
rect 0 1484 364 1512
rect 532 1484 672 1512
rect 784 1484 1568 1512
rect 1792 1540 3024 1568
rect 3192 1540 3584 1568
rect 1792 1512 2548 1540
rect 2660 1512 3024 1540
rect 1792 1484 2492 1512
rect 2660 1484 2744 1512
rect 0 1456 392 1484
rect 532 1456 644 1484
rect 812 1456 2464 1484
rect 2660 1456 2716 1484
rect 2856 1456 3024 1512
rect 3164 1484 3584 1540
rect 3192 1456 3584 1484
rect 0 1428 420 1456
rect 532 1428 588 1456
rect 812 1428 924 1456
rect 1008 1428 2436 1456
rect 2856 1428 3052 1456
rect 3220 1428 3584 1456
rect 0 1372 392 1428
rect 532 1400 560 1428
rect 840 1400 896 1428
rect 0 1316 364 1372
rect 504 1344 560 1400
rect 700 1372 728 1400
rect 672 1344 728 1372
rect 1008 1372 2408 1428
rect 2828 1400 3080 1428
rect 2548 1372 2576 1400
rect 2800 1372 3108 1400
rect 3248 1372 3584 1428
rect 1008 1344 2072 1372
rect 2156 1344 2408 1372
rect 2520 1344 2576 1372
rect 2744 1344 3136 1372
rect 3276 1344 3584 1372
rect 0 1064 336 1316
rect 476 1288 756 1344
rect 980 1316 1708 1344
rect 1792 1316 2016 1344
rect 924 1288 1680 1316
rect 1820 1288 1988 1316
rect 2156 1288 2576 1344
rect 2716 1316 3164 1344
rect 2688 1288 3164 1316
rect 3304 1288 3584 1344
rect 448 1260 1652 1288
rect 2156 1260 3192 1288
rect 448 1232 1400 1260
rect 1540 1232 1596 1260
rect 2100 1232 3192 1260
rect 420 1176 1400 1232
rect 2072 1204 3136 1232
rect 3332 1204 3584 1288
rect 1736 1176 1820 1204
rect 1988 1176 2688 1204
rect 2800 1176 3080 1204
rect 3304 1176 3584 1204
rect 420 1148 1456 1176
rect 1680 1148 2660 1176
rect 2800 1148 2912 1176
rect 3276 1148 3584 1176
rect 504 1120 644 1148
rect 868 1120 2632 1148
rect 3220 1120 3584 1148
rect 924 1092 2576 1120
rect 2772 1092 2800 1120
rect 3136 1092 3584 1120
rect 952 1064 2520 1092
rect 2744 1064 2800 1092
rect 2996 1064 3584 1092
rect 0 1036 420 1064
rect 728 1036 784 1064
rect 1008 1036 2464 1064
rect 2716 1036 3584 1064
rect 0 1008 840 1036
rect 1064 1008 2380 1036
rect 2660 1008 3584 1036
rect 0 980 868 1008
rect 1288 980 2296 1008
rect 2604 980 3584 1008
rect 0 952 924 980
rect 1344 952 2296 980
rect 2520 952 3584 980
rect 0 924 980 952
rect 1512 924 2296 952
rect 2436 924 3584 952
rect 0 868 1036 924
rect 1148 896 1204 924
rect 1512 896 3584 924
rect 1176 868 1288 896
rect 1512 868 2408 896
rect 0 812 1064 868
rect 1176 840 2408 868
rect 2520 840 3584 896
rect 1204 812 2408 840
rect 2548 812 3584 840
rect 0 756 1092 812
rect 1232 784 2436 812
rect 1260 756 2436 784
rect 0 728 1120 756
rect 1288 728 2464 756
rect 2576 728 3584 812
rect 0 700 1148 728
rect 0 672 1176 700
rect 1316 672 2492 728
rect 2604 672 3584 728
rect 0 644 1204 672
rect 0 588 1176 644
rect 1316 588 2520 672
rect 0 560 1148 588
rect 1288 560 2548 588
rect 2632 560 3584 672
rect 0 532 1120 560
rect 1260 532 2548 560
rect 0 504 1092 532
rect 0 392 1064 504
rect 1232 476 2548 532
rect 2660 476 3584 560
rect 1372 448 2576 476
rect 1400 392 2576 448
rect 0 308 1260 392
rect 1400 364 2604 392
rect 2688 364 3584 476
rect 1372 308 2604 364
rect 0 224 1232 308
rect 1344 252 2632 308
rect 2716 252 3584 364
rect 0 28 1204 224
rect 1316 168 2632 252
rect 1288 28 2660 168
rect 2744 28 3584 252
rect 0 0 3584 28
<< obsm3 >>
rect 0 0 3584 3584
<< obsm4 >>
rect 0 0 3584 3584
<< obsm5 >>
rect 0 0 3584 3584
<< properties >>
string FIXED_BBOX 0 0 3584 3584
<< end >>
