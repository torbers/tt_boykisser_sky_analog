VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO my_logo
  CLASS BLOCK ;
  FOREIGN my_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.840 BY 35.840 ;
  OBS
      LAYER met1 ;
        RECT 0.000 35.560 35.840 35.840 ;
        RECT 0.000 35.280 29.960 35.560 ;
      LAYER met1 ;
        RECT 29.960 35.280 31.360 35.560 ;
      LAYER met1 ;
        RECT 0.000 34.160 4.200 35.280 ;
      LAYER met1 ;
        RECT 4.200 35.000 5.600 35.280 ;
      LAYER met1 ;
        RECT 5.600 35.000 29.120 35.280 ;
      LAYER met1 ;
        RECT 29.120 35.000 31.360 35.280 ;
      LAYER met1 ;
        RECT 31.360 35.000 35.840 35.560 ;
      LAYER met1 ;
        RECT 4.200 34.720 6.720 35.000 ;
      LAYER met1 ;
        RECT 6.720 34.720 28.560 35.000 ;
      LAYER met1 ;
        RECT 28.560 34.720 31.640 35.000 ;
        RECT 4.200 34.440 7.560 34.720 ;
      LAYER met1 ;
        RECT 7.560 34.440 27.720 34.720 ;
      LAYER met1 ;
        RECT 27.720 34.440 31.640 34.720 ;
        RECT 4.200 34.160 8.120 34.440 ;
      LAYER met1 ;
        RECT 8.120 34.160 27.160 34.440 ;
      LAYER met1 ;
        RECT 27.160 34.160 29.960 34.440 ;
      LAYER met1 ;
        RECT 29.960 34.160 30.800 34.440 ;
      LAYER met1 ;
        RECT 30.800 34.160 31.640 34.440 ;
      LAYER met1 ;
        RECT 31.640 34.160 35.840 35.000 ;
        RECT 0.000 33.040 3.920 34.160 ;
      LAYER met1 ;
        RECT 3.920 33.320 5.040 34.160 ;
      LAYER met1 ;
        RECT 5.040 33.880 6.160 34.160 ;
      LAYER met1 ;
        RECT 6.160 33.880 8.400 34.160 ;
      LAYER met1 ;
        RECT 8.400 33.880 26.600 34.160 ;
      LAYER met1 ;
        RECT 26.600 33.880 29.120 34.160 ;
      LAYER met1 ;
        RECT 29.120 33.880 30.800 34.160 ;
        RECT 5.040 33.600 6.720 33.880 ;
      LAYER met1 ;
        RECT 6.720 33.600 8.680 33.880 ;
      LAYER met1 ;
        RECT 8.680 33.600 26.040 33.880 ;
      LAYER met1 ;
        RECT 26.040 33.600 28.560 33.880 ;
      LAYER met1 ;
        RECT 28.560 33.600 30.800 33.880 ;
      LAYER met1 ;
        RECT 30.800 33.600 31.920 34.160 ;
      LAYER met1 ;
        RECT 5.040 33.320 7.280 33.600 ;
      LAYER met1 ;
        RECT 7.280 33.320 8.960 33.600 ;
      LAYER met1 ;
        RECT 8.960 33.320 25.760 33.600 ;
      LAYER met1 ;
        RECT 25.760 33.320 28.000 33.600 ;
      LAYER met1 ;
        RECT 28.000 33.320 31.080 33.600 ;
      LAYER met1 ;
        RECT 31.080 33.320 31.920 33.600 ;
      LAYER met1 ;
        RECT 31.920 33.320 35.840 34.160 ;
      LAYER met1 ;
        RECT 3.920 33.040 4.760 33.320 ;
      LAYER met1 ;
        RECT 4.760 33.040 7.560 33.320 ;
      LAYER met1 ;
        RECT 7.560 33.040 9.240 33.320 ;
      LAYER met1 ;
        RECT 9.240 33.040 13.720 33.320 ;
      LAYER met1 ;
        RECT 13.720 33.040 14.560 33.320 ;
      LAYER met1 ;
        RECT 14.560 33.040 25.200 33.320 ;
      LAYER met1 ;
        RECT 25.200 33.040 27.440 33.320 ;
      LAYER met1 ;
        RECT 27.440 33.040 31.080 33.320 ;
        RECT 0.000 31.640 3.640 33.040 ;
      LAYER met1 ;
        RECT 3.640 32.480 4.760 33.040 ;
      LAYER met1 ;
        RECT 4.760 32.760 7.840 33.040 ;
      LAYER met1 ;
        RECT 7.840 32.760 9.800 33.040 ;
      LAYER met1 ;
        RECT 9.800 32.760 13.720 33.040 ;
      LAYER met1 ;
        RECT 13.720 32.760 16.800 33.040 ;
      LAYER met1 ;
        RECT 16.800 32.760 24.920 33.040 ;
      LAYER met1 ;
        RECT 24.920 32.760 26.880 33.040 ;
      LAYER met1 ;
        RECT 26.880 32.760 31.080 33.040 ;
      LAYER met1 ;
        RECT 31.080 32.760 32.200 33.320 ;
      LAYER met1 ;
        RECT 4.760 32.480 8.400 32.760 ;
      LAYER met1 ;
        RECT 8.400 32.480 10.080 32.760 ;
      LAYER met1 ;
        RECT 10.080 32.480 13.720 32.760 ;
      LAYER met1 ;
        RECT 13.720 32.480 17.640 32.760 ;
      LAYER met1 ;
        RECT 17.640 32.480 24.640 32.760 ;
      LAYER met1 ;
        RECT 24.640 32.480 26.320 32.760 ;
      LAYER met1 ;
        RECT 26.320 32.480 31.360 32.760 ;
      LAYER met1 ;
        RECT 31.360 32.480 32.200 32.760 ;
      LAYER met1 ;
        RECT 32.200 32.480 35.840 33.320 ;
      LAYER met1 ;
        RECT 3.640 31.640 4.480 32.480 ;
      LAYER met1 ;
        RECT 4.480 32.200 8.680 32.480 ;
      LAYER met1 ;
        RECT 8.680 32.200 10.640 32.480 ;
      LAYER met1 ;
        RECT 10.640 32.200 13.720 32.480 ;
      LAYER met1 ;
        RECT 13.720 32.200 18.480 32.480 ;
      LAYER met1 ;
        RECT 18.480 32.200 24.080 32.480 ;
      LAYER met1 ;
        RECT 24.080 32.200 26.040 32.480 ;
      LAYER met1 ;
        RECT 26.040 32.200 31.360 32.480 ;
        RECT 4.480 31.920 8.960 32.200 ;
      LAYER met1 ;
        RECT 8.960 31.920 10.920 32.200 ;
      LAYER met1 ;
        RECT 10.920 31.920 13.720 32.200 ;
      LAYER met1 ;
        RECT 13.720 31.920 14.840 32.200 ;
      LAYER met1 ;
        RECT 14.840 31.920 15.960 32.200 ;
      LAYER met1 ;
        RECT 15.960 31.920 19.320 32.200 ;
      LAYER met1 ;
        RECT 19.320 31.920 23.800 32.200 ;
      LAYER met1 ;
        RECT 23.800 31.920 25.760 32.200 ;
      LAYER met1 ;
        RECT 25.760 31.920 31.360 32.200 ;
        RECT 4.480 31.640 9.520 31.920 ;
      LAYER met1 ;
        RECT 9.520 31.640 11.200 31.920 ;
      LAYER met1 ;
        RECT 11.200 31.640 14.000 31.920 ;
      LAYER met1 ;
        RECT 14.000 31.640 14.840 31.920 ;
      LAYER met1 ;
        RECT 14.840 31.640 17.080 31.920 ;
      LAYER met1 ;
        RECT 17.080 31.640 19.880 31.920 ;
      LAYER met1 ;
        RECT 19.880 31.640 23.800 31.920 ;
      LAYER met1 ;
        RECT 23.800 31.640 25.480 31.920 ;
      LAYER met1 ;
        RECT 25.480 31.640 31.360 31.920 ;
      LAYER met1 ;
        RECT 31.360 31.640 32.480 32.480 ;
      LAYER met1 ;
        RECT 0.000 30.240 3.360 31.640 ;
      LAYER met1 ;
        RECT 3.360 31.080 4.480 31.640 ;
      LAYER met1 ;
        RECT 4.480 31.360 9.800 31.640 ;
      LAYER met1 ;
        RECT 9.800 31.360 11.480 31.640 ;
      LAYER met1 ;
        RECT 11.480 31.360 14.000 31.640 ;
        RECT 4.480 31.080 10.080 31.360 ;
      LAYER met1 ;
        RECT 10.080 31.080 11.760 31.360 ;
      LAYER met1 ;
        RECT 11.760 31.080 14.000 31.360 ;
      LAYER met1 ;
        RECT 14.000 31.080 15.120 31.640 ;
      LAYER met1 ;
        RECT 15.120 31.360 17.920 31.640 ;
      LAYER met1 ;
        RECT 17.920 31.360 20.440 31.640 ;
      LAYER met1 ;
        RECT 20.440 31.360 23.520 31.640 ;
      LAYER met1 ;
        RECT 23.520 31.360 25.200 31.640 ;
      LAYER met1 ;
        RECT 25.200 31.360 31.640 31.640 ;
      LAYER met1 ;
        RECT 31.640 31.360 32.480 31.640 ;
      LAYER met1 ;
        RECT 32.480 31.360 35.840 32.480 ;
        RECT 15.120 31.080 18.480 31.360 ;
      LAYER met1 ;
        RECT 18.480 31.080 21.000 31.360 ;
      LAYER met1 ;
        RECT 21.000 31.080 23.520 31.360 ;
      LAYER met1 ;
        RECT 23.520 31.080 24.920 31.360 ;
      LAYER met1 ;
        RECT 24.920 31.080 31.640 31.360 ;
      LAYER met1 ;
        RECT 3.360 30.240 4.200 31.080 ;
      LAYER met1 ;
        RECT 4.200 30.800 10.360 31.080 ;
      LAYER met1 ;
        RECT 10.360 30.800 12.040 31.080 ;
      LAYER met1 ;
        RECT 4.200 30.520 10.640 30.800 ;
      LAYER met1 ;
        RECT 10.640 30.520 12.040 30.800 ;
      LAYER met1 ;
        RECT 12.040 30.520 14.280 31.080 ;
      LAYER met1 ;
        RECT 14.280 30.520 15.400 31.080 ;
      LAYER met1 ;
        RECT 15.400 30.800 19.040 31.080 ;
      LAYER met1 ;
        RECT 19.040 30.800 21.280 31.080 ;
      LAYER met1 ;
        RECT 21.280 30.800 23.240 31.080 ;
      LAYER met1 ;
        RECT 23.240 30.800 24.360 31.080 ;
      LAYER met1 ;
        RECT 15.400 30.520 19.600 30.800 ;
      LAYER met1 ;
        RECT 19.600 30.520 21.560 30.800 ;
      LAYER met1 ;
        RECT 21.560 30.520 22.960 30.800 ;
      LAYER met1 ;
        RECT 22.960 30.520 24.360 30.800 ;
      LAYER met1 ;
        RECT 24.360 30.520 31.640 31.080 ;
      LAYER met1 ;
        RECT 31.640 30.520 32.760 31.360 ;
      LAYER met1 ;
        RECT 4.200 30.240 10.920 30.520 ;
      LAYER met1 ;
        RECT 10.920 30.240 12.320 30.520 ;
      LAYER met1 ;
        RECT 12.320 30.240 14.280 30.520 ;
      LAYER met1 ;
        RECT 14.280 30.240 15.680 30.520 ;
      LAYER met1 ;
        RECT 15.680 30.240 20.160 30.520 ;
      LAYER met1 ;
        RECT 20.160 30.240 21.840 30.520 ;
      LAYER met1 ;
        RECT 21.840 30.240 22.960 30.520 ;
      LAYER met1 ;
        RECT 22.960 30.240 24.080 30.520 ;
      LAYER met1 ;
        RECT 0.000 28.000 3.080 30.240 ;
      LAYER met1 ;
        RECT 3.080 29.680 4.200 30.240 ;
      LAYER met1 ;
        RECT 4.200 29.960 11.200 30.240 ;
      LAYER met1 ;
        RECT 11.200 29.960 12.600 30.240 ;
      LAYER met1 ;
        RECT 12.600 29.960 14.560 30.240 ;
      LAYER met1 ;
        RECT 14.560 29.960 15.960 30.240 ;
      LAYER met1 ;
        RECT 15.960 29.960 20.440 30.240 ;
      LAYER met1 ;
        RECT 20.440 29.960 22.400 30.240 ;
      LAYER met1 ;
        RECT 22.400 29.960 22.680 30.240 ;
      LAYER met1 ;
        RECT 22.680 29.960 24.080 30.240 ;
      LAYER met1 ;
        RECT 24.080 29.960 31.920 30.520 ;
      LAYER met1 ;
        RECT 31.920 29.960 32.760 30.520 ;
      LAYER met1 ;
        RECT 32.760 29.960 35.840 31.360 ;
        RECT 4.200 29.680 11.480 29.960 ;
      LAYER met1 ;
        RECT 11.480 29.680 12.880 29.960 ;
      LAYER met1 ;
        RECT 12.880 29.680 14.560 29.960 ;
      LAYER met1 ;
        RECT 14.560 29.680 16.240 29.960 ;
      LAYER met1 ;
        RECT 16.240 29.680 21.000 29.960 ;
      LAYER met1 ;
        RECT 21.000 29.680 23.800 29.960 ;
        RECT 3.080 28.000 3.920 29.680 ;
      LAYER met1 ;
        RECT 3.920 29.400 11.760 29.680 ;
      LAYER met1 ;
        RECT 11.760 29.400 13.160 29.680 ;
      LAYER met1 ;
        RECT 13.160 29.400 14.840 29.680 ;
      LAYER met1 ;
        RECT 14.840 29.400 16.520 29.680 ;
      LAYER met1 ;
        RECT 16.520 29.400 21.280 29.680 ;
      LAYER met1 ;
        RECT 21.280 29.400 23.800 29.680 ;
      LAYER met1 ;
        RECT 23.800 29.400 31.920 29.960 ;
      LAYER met1 ;
        RECT 31.920 29.400 33.040 29.960 ;
      LAYER met1 ;
        RECT 3.920 29.120 12.040 29.400 ;
      LAYER met1 ;
        RECT 12.040 29.120 13.440 29.400 ;
      LAYER met1 ;
        RECT 13.440 29.120 15.120 29.400 ;
      LAYER met1 ;
        RECT 15.120 29.120 16.520 29.400 ;
      LAYER met1 ;
        RECT 16.520 29.120 21.560 29.400 ;
      LAYER met1 ;
        RECT 21.560 29.120 23.520 29.400 ;
      LAYER met1 ;
        RECT 3.920 28.560 12.320 29.120 ;
      LAYER met1 ;
        RECT 12.320 28.840 13.720 29.120 ;
      LAYER met1 ;
        RECT 13.720 28.840 15.400 29.120 ;
      LAYER met1 ;
        RECT 15.400 28.840 16.800 29.120 ;
      LAYER met1 ;
        RECT 16.800 28.840 21.840 29.120 ;
      LAYER met1 ;
        RECT 21.840 28.840 23.520 29.120 ;
      LAYER met1 ;
        RECT 23.520 28.840 32.200 29.400 ;
      LAYER met1 ;
        RECT 32.200 28.840 33.040 29.400 ;
      LAYER met1 ;
        RECT 33.040 28.840 35.840 29.960 ;
      LAYER met1 ;
        RECT 12.320 28.560 14.000 28.840 ;
      LAYER met1 ;
        RECT 14.000 28.560 14.560 28.840 ;
      LAYER met1 ;
        RECT 14.560 28.560 16.800 28.840 ;
      LAYER met1 ;
        RECT 16.800 28.560 22.120 28.840 ;
      LAYER met1 ;
        RECT 22.120 28.560 23.240 28.840 ;
      LAYER met1 ;
        RECT 3.920 28.280 12.600 28.560 ;
      LAYER met1 ;
        RECT 12.600 28.280 16.800 28.560 ;
      LAYER met1 ;
        RECT 16.800 28.280 22.400 28.560 ;
        RECT 3.920 28.000 12.880 28.280 ;
      LAYER met1 ;
        RECT 12.880 28.000 16.240 28.280 ;
      LAYER met1 ;
        RECT 16.240 28.000 22.400 28.280 ;
      LAYER met1 ;
        RECT 22.400 28.000 23.240 28.560 ;
      LAYER met1 ;
        RECT 23.240 28.000 32.200 28.840 ;
      LAYER met1 ;
        RECT 32.200 28.000 33.320 28.840 ;
      LAYER met1 ;
        RECT 0.000 26.320 2.800 28.000 ;
      LAYER met1 ;
        RECT 2.800 27.440 3.920 28.000 ;
      LAYER met1 ;
        RECT 3.920 27.720 13.440 28.000 ;
      LAYER met1 ;
        RECT 13.440 27.720 15.120 28.000 ;
      LAYER met1 ;
        RECT 15.120 27.720 32.480 28.000 ;
        RECT 3.920 27.440 13.160 27.720 ;
      LAYER met1 ;
        RECT 13.160 27.440 14.840 27.720 ;
      LAYER met1 ;
        RECT 14.840 27.440 32.480 27.720 ;
      LAYER met1 ;
        RECT 2.800 26.320 3.640 27.440 ;
      LAYER met1 ;
        RECT 3.640 27.160 12.880 27.440 ;
      LAYER met1 ;
        RECT 12.880 27.160 14.560 27.440 ;
      LAYER met1 ;
        RECT 14.560 27.160 32.480 27.440 ;
      LAYER met1 ;
        RECT 32.480 27.160 33.320 28.000 ;
      LAYER met1 ;
        RECT 33.320 27.160 35.840 28.840 ;
        RECT 0.000 23.800 2.520 26.320 ;
      LAYER met1 ;
        RECT 2.520 25.480 3.640 26.320 ;
      LAYER met1 ;
        RECT 3.640 26.040 12.600 27.160 ;
      LAYER met1 ;
        RECT 12.600 26.880 14.280 27.160 ;
      LAYER met1 ;
        RECT 14.280 26.880 32.480 27.160 ;
      LAYER met1 ;
        RECT 12.600 26.600 17.360 26.880 ;
      LAYER met1 ;
        RECT 17.360 26.600 32.480 26.880 ;
      LAYER met1 ;
        RECT 32.480 26.600 33.600 27.160 ;
        RECT 12.600 26.040 18.200 26.600 ;
      LAYER met1 ;
        RECT 3.640 25.760 16.520 26.040 ;
      LAYER met1 ;
        RECT 16.520 25.760 18.200 26.040 ;
      LAYER met1 ;
        RECT 18.200 25.760 32.760 26.600 ;
      LAYER met1 ;
        RECT 32.760 26.320 33.600 26.600 ;
      LAYER met1 ;
        RECT 33.600 26.320 35.840 27.160 ;
        RECT 3.640 25.480 32.760 25.760 ;
      LAYER met1 ;
        RECT 32.760 25.480 33.880 26.320 ;
      LAYER met1 ;
        RECT 33.880 25.480 35.840 26.320 ;
      LAYER met1 ;
        RECT 2.520 24.640 3.360 25.480 ;
      LAYER met1 ;
        RECT 3.360 24.640 32.760 25.480 ;
      LAYER met1 ;
        RECT 2.520 23.800 3.640 24.640 ;
      LAYER met1 ;
        RECT 3.640 24.360 32.760 24.640 ;
      LAYER met1 ;
        RECT 32.760 24.360 33.600 25.480 ;
      LAYER met1 ;
        RECT 0.000 22.680 2.800 23.800 ;
      LAYER met1 ;
        RECT 2.800 23.520 3.640 23.800 ;
      LAYER met1 ;
        RECT 3.640 23.520 32.480 24.360 ;
      LAYER met1 ;
        RECT 32.480 23.520 33.600 24.360 ;
      LAYER met1 ;
        RECT 33.600 23.520 35.840 25.480 ;
      LAYER met1 ;
        RECT 2.800 22.680 3.920 23.520 ;
      LAYER met1 ;
        RECT 3.920 22.960 32.480 23.520 ;
      LAYER met1 ;
        RECT 32.480 22.960 33.320 23.520 ;
      LAYER met1 ;
        RECT 3.920 22.680 32.200 22.960 ;
        RECT 0.000 21.840 3.080 22.680 ;
      LAYER met1 ;
        RECT 3.080 22.120 4.200 22.680 ;
      LAYER met1 ;
        RECT 4.200 22.400 32.200 22.680 ;
      LAYER met1 ;
        RECT 32.200 22.400 33.320 22.960 ;
      LAYER met1 ;
        RECT 33.320 22.400 35.840 23.520 ;
        RECT 4.200 22.120 31.920 22.400 ;
      LAYER met1 ;
        RECT 31.920 22.120 33.040 22.400 ;
        RECT 3.080 21.840 4.480 22.120 ;
      LAYER met1 ;
        RECT 4.480 21.840 31.640 22.120 ;
      LAYER met1 ;
        RECT 31.640 21.840 33.040 22.120 ;
      LAYER met1 ;
        RECT 33.040 21.840 35.840 22.400 ;
        RECT 0.000 21.280 3.360 21.840 ;
      LAYER met1 ;
        RECT 3.360 21.280 4.480 21.840 ;
      LAYER met1 ;
        RECT 4.480 21.560 22.120 21.840 ;
      LAYER met1 ;
        RECT 22.120 21.560 28.000 21.840 ;
      LAYER met1 ;
        RECT 28.000 21.560 31.640 21.840 ;
      LAYER met1 ;
        RECT 31.640 21.560 32.760 21.840 ;
      LAYER met1 ;
        RECT 4.480 21.280 21.560 21.560 ;
      LAYER met1 ;
        RECT 21.560 21.280 28.000 21.560 ;
      LAYER met1 ;
        RECT 28.000 21.280 31.360 21.560 ;
      LAYER met1 ;
        RECT 31.360 21.280 32.760 21.560 ;
      LAYER met1 ;
        RECT 32.760 21.280 35.840 21.840 ;
        RECT 0.000 20.440 3.640 21.280 ;
      LAYER met1 ;
        RECT 3.640 20.440 4.760 21.280 ;
      LAYER met1 ;
        RECT 4.760 20.440 7.560 21.280 ;
      LAYER met1 ;
        RECT 7.560 21.000 14.280 21.280 ;
      LAYER met1 ;
        RECT 14.280 21.000 21.000 21.280 ;
      LAYER met1 ;
        RECT 21.000 21.000 28.000 21.280 ;
      LAYER met1 ;
        RECT 28.000 21.000 31.080 21.280 ;
      LAYER met1 ;
        RECT 31.080 21.000 32.480 21.280 ;
        RECT 7.560 20.440 14.840 21.000 ;
      LAYER met1 ;
        RECT 14.840 20.440 21.000 21.000 ;
      LAYER met1 ;
        RECT 21.000 20.440 24.360 21.000 ;
      LAYER met1 ;
        RECT 24.360 20.440 25.760 21.000 ;
      LAYER met1 ;
        RECT 25.760 20.440 27.160 21.000 ;
      LAYER met1 ;
        RECT 27.160 20.720 30.800 21.000 ;
      LAYER met1 ;
        RECT 30.800 20.720 32.480 21.000 ;
      LAYER met1 ;
        RECT 32.480 20.720 35.840 21.280 ;
        RECT 27.160 20.440 30.520 20.720 ;
      LAYER met1 ;
        RECT 30.520 20.440 32.200 20.720 ;
      LAYER met1 ;
        RECT 32.200 20.440 35.840 20.720 ;
        RECT 0.000 19.880 3.920 20.440 ;
      LAYER met1 ;
        RECT 3.920 19.880 5.040 20.440 ;
      LAYER met1 ;
        RECT 5.040 20.160 8.400 20.440 ;
      LAYER met1 ;
        RECT 8.400 20.160 9.800 20.440 ;
      LAYER met1 ;
        RECT 5.040 19.880 8.120 20.160 ;
      LAYER met1 ;
        RECT 8.120 19.880 9.800 20.160 ;
      LAYER met1 ;
        RECT 9.800 19.880 11.200 20.440 ;
        RECT 0.000 19.040 4.200 19.880 ;
      LAYER met1 ;
        RECT 4.200 19.320 5.320 19.880 ;
      LAYER met1 ;
        RECT 5.320 19.600 8.120 19.880 ;
      LAYER met1 ;
        RECT 8.120 19.600 9.520 19.880 ;
      LAYER met1 ;
        RECT 9.520 19.600 11.200 19.880 ;
        RECT 5.320 19.320 7.840 19.600 ;
      LAYER met1 ;
        RECT 7.840 19.320 9.240 19.600 ;
      LAYER met1 ;
        RECT 9.240 19.320 11.200 19.600 ;
      LAYER met1 ;
        RECT 4.200 19.040 5.600 19.320 ;
      LAYER met1 ;
        RECT 0.000 18.760 4.480 19.040 ;
      LAYER met1 ;
        RECT 4.480 18.760 5.600 19.040 ;
      LAYER met1 ;
        RECT 5.600 18.760 7.840 19.320 ;
      LAYER met1 ;
        RECT 7.840 18.760 8.960 19.320 ;
      LAYER met1 ;
        RECT 8.960 18.760 11.200 19.320 ;
        RECT 0.000 17.360 1.680 18.760 ;
      LAYER met1 ;
        RECT 1.680 18.480 2.520 18.760 ;
      LAYER met1 ;
        RECT 2.520 18.480 4.480 18.760 ;
      LAYER met1 ;
        RECT 4.480 18.480 5.880 18.760 ;
        RECT 1.680 18.200 3.360 18.480 ;
      LAYER met1 ;
        RECT 3.360 18.200 4.760 18.480 ;
      LAYER met1 ;
        RECT 4.760 18.200 5.880 18.480 ;
      LAYER met1 ;
        RECT 5.880 18.200 7.560 18.760 ;
      LAYER met1 ;
        RECT 1.680 17.360 7.000 18.200 ;
      LAYER met1 ;
        RECT 7.000 17.360 7.560 18.200 ;
      LAYER met1 ;
        RECT 7.560 17.920 8.680 18.760 ;
      LAYER met1 ;
        RECT 8.680 17.920 11.200 18.760 ;
      LAYER met1 ;
        RECT 11.200 17.920 15.120 20.440 ;
      LAYER met1 ;
        RECT 15.120 17.920 20.720 20.440 ;
        RECT 0.000 16.800 1.960 17.360 ;
      LAYER met1 ;
        RECT 1.960 17.080 3.080 17.360 ;
      LAYER met1 ;
        RECT 3.080 17.080 7.560 17.360 ;
      LAYER met1 ;
        RECT 7.560 17.080 8.400 17.920 ;
      LAYER met1 ;
        RECT 8.400 17.080 11.200 17.920 ;
      LAYER met1 ;
        RECT 11.200 17.080 14.840 17.920 ;
      LAYER met1 ;
        RECT 14.840 17.080 20.720 17.920 ;
      LAYER met1 ;
        RECT 20.720 17.080 24.360 20.440 ;
      LAYER met1 ;
        RECT 24.360 20.160 26.040 20.440 ;
      LAYER met1 ;
        RECT 26.040 20.160 27.160 20.440 ;
      LAYER met1 ;
        RECT 27.160 20.160 30.240 20.440 ;
      LAYER met1 ;
        RECT 30.240 20.160 31.920 20.440 ;
      LAYER met1 ;
        RECT 31.920 20.160 35.840 20.440 ;
        RECT 24.360 19.600 26.320 20.160 ;
      LAYER met1 ;
        RECT 26.320 19.600 27.440 20.160 ;
      LAYER met1 ;
        RECT 27.440 19.880 30.240 20.160 ;
      LAYER met1 ;
        RECT 30.240 19.880 31.640 20.160 ;
      LAYER met1 ;
        RECT 31.640 19.880 35.840 20.160 ;
        RECT 27.440 19.600 29.680 19.880 ;
      LAYER met1 ;
        RECT 29.680 19.600 31.360 19.880 ;
      LAYER met1 ;
        RECT 31.360 19.600 35.840 19.880 ;
        RECT 24.360 18.200 26.600 19.600 ;
      LAYER met1 ;
        RECT 26.600 19.040 27.440 19.600 ;
      LAYER met1 ;
        RECT 27.440 19.320 29.400 19.600 ;
      LAYER met1 ;
        RECT 29.400 19.320 34.440 19.600 ;
      LAYER met1 ;
        RECT 27.440 19.040 29.120 19.320 ;
      LAYER met1 ;
        RECT 26.600 18.200 27.720 19.040 ;
      LAYER met1 ;
        RECT 27.720 18.200 29.120 19.040 ;
      LAYER met1 ;
        RECT 29.120 18.760 34.440 19.320 ;
        RECT 29.120 18.480 31.920 18.760 ;
      LAYER met1 ;
        RECT 31.920 18.480 33.040 18.760 ;
      LAYER met1 ;
        RECT 33.040 18.480 34.440 18.760 ;
      LAYER met1 ;
        RECT 34.440 18.480 35.840 19.600 ;
      LAYER met1 ;
        RECT 29.120 18.200 29.960 18.480 ;
      LAYER met1 ;
        RECT 29.960 18.200 32.760 18.480 ;
      LAYER met1 ;
        RECT 32.760 18.200 34.160 18.480 ;
      LAYER met1 ;
        RECT 34.160 18.200 35.840 18.480 ;
        RECT 24.360 17.360 26.880 18.200 ;
      LAYER met1 ;
        RECT 26.880 17.360 27.720 18.200 ;
      LAYER met1 ;
        RECT 27.720 17.920 32.760 18.200 ;
      LAYER met1 ;
        RECT 32.760 17.920 33.880 18.200 ;
      LAYER met1 ;
        RECT 27.720 17.640 32.480 17.920 ;
      LAYER met1 ;
        RECT 32.480 17.640 33.880 17.920 ;
      LAYER met1 ;
        RECT 33.880 17.640 35.840 18.200 ;
        RECT 27.720 17.360 32.200 17.640 ;
      LAYER met1 ;
        RECT 32.200 17.360 33.600 17.640 ;
      LAYER met1 ;
        RECT 33.600 17.360 35.840 17.640 ;
        RECT 24.360 17.080 26.600 17.360 ;
      LAYER met1 ;
        RECT 1.960 16.800 3.360 17.080 ;
      LAYER met1 ;
        RECT 3.360 16.800 7.560 17.080 ;
        RECT 0.000 16.520 2.240 16.800 ;
      LAYER met1 ;
        RECT 2.240 16.520 3.640 16.800 ;
      LAYER met1 ;
        RECT 3.640 16.520 7.560 16.800 ;
        RECT 0.000 15.960 2.520 16.520 ;
      LAYER met1 ;
        RECT 2.520 16.240 3.920 16.520 ;
      LAYER met1 ;
        RECT 3.920 16.240 7.560 16.520 ;
      LAYER met1 ;
        RECT 7.560 16.240 8.680 17.080 ;
      LAYER met1 ;
        RECT 8.680 16.520 11.480 17.080 ;
      LAYER met1 ;
        RECT 11.480 16.520 14.560 17.080 ;
      LAYER met1 ;
        RECT 14.560 16.520 21.000 17.080 ;
      LAYER met1 ;
        RECT 21.000 16.520 24.080 17.080 ;
      LAYER met1 ;
        RECT 24.080 16.520 26.600 17.080 ;
      LAYER met1 ;
        RECT 26.600 16.520 27.720 17.360 ;
      LAYER met1 ;
        RECT 27.720 17.080 31.920 17.360 ;
      LAYER met1 ;
        RECT 31.920 17.080 33.320 17.360 ;
      LAYER met1 ;
        RECT 33.320 17.080 35.840 17.360 ;
        RECT 27.720 16.800 31.640 17.080 ;
      LAYER met1 ;
        RECT 31.640 16.800 33.040 17.080 ;
      LAYER met1 ;
        RECT 33.040 16.800 35.840 17.080 ;
        RECT 27.720 16.520 31.360 16.800 ;
      LAYER met1 ;
        RECT 31.360 16.520 32.760 16.800 ;
      LAYER met1 ;
        RECT 8.680 16.240 11.760 16.520 ;
      LAYER met1 ;
        RECT 11.760 16.240 14.280 16.520 ;
      LAYER met1 ;
        RECT 14.280 16.240 21.280 16.520 ;
      LAYER met1 ;
        RECT 21.280 16.240 23.800 16.520 ;
      LAYER met1 ;
        RECT 23.800 16.240 26.600 16.520 ;
      LAYER met1 ;
        RECT 2.520 15.960 4.200 16.240 ;
      LAYER met1 ;
        RECT 4.200 15.960 7.840 16.240 ;
        RECT 0.000 15.680 2.800 15.960 ;
      LAYER met1 ;
        RECT 2.800 15.680 4.480 15.960 ;
      LAYER met1 ;
        RECT 4.480 15.680 7.840 15.960 ;
        RECT 0.000 15.400 3.080 15.680 ;
      LAYER met1 ;
        RECT 3.080 15.400 4.760 15.680 ;
      LAYER met1 ;
        RECT 4.760 15.400 7.840 15.680 ;
      LAYER met1 ;
        RECT 7.840 15.400 8.960 16.240 ;
      LAYER met1 ;
        RECT 8.960 15.960 11.760 16.240 ;
      LAYER met1 ;
        RECT 11.760 15.960 14.000 16.240 ;
      LAYER met1 ;
        RECT 14.000 15.960 21.840 16.240 ;
      LAYER met1 ;
        RECT 21.840 15.960 23.240 16.240 ;
      LAYER met1 ;
        RECT 23.240 15.960 26.600 16.240 ;
      LAYER met1 ;
        RECT 26.600 15.960 27.440 16.520 ;
      LAYER met1 ;
        RECT 27.440 16.240 31.080 16.520 ;
      LAYER met1 ;
        RECT 31.080 16.240 32.760 16.520 ;
      LAYER met1 ;
        RECT 32.760 16.240 35.840 16.800 ;
        RECT 27.440 15.960 30.800 16.240 ;
      LAYER met1 ;
        RECT 30.800 15.960 32.480 16.240 ;
      LAYER met1 ;
        RECT 32.480 15.960 35.840 16.240 ;
        RECT 8.960 15.680 12.040 15.960 ;
      LAYER met1 ;
        RECT 12.040 15.680 13.720 15.960 ;
      LAYER met1 ;
        RECT 13.720 15.680 30.520 15.960 ;
      LAYER met1 ;
        RECT 30.520 15.680 32.200 15.960 ;
      LAYER met1 ;
        RECT 32.200 15.680 35.840 15.960 ;
        RECT 0.000 15.120 3.360 15.400 ;
      LAYER met1 ;
        RECT 3.360 15.120 5.040 15.400 ;
      LAYER met1 ;
        RECT 5.040 15.120 8.120 15.400 ;
      LAYER met1 ;
        RECT 8.120 15.120 8.960 15.400 ;
      LAYER met1 ;
        RECT 8.960 15.120 15.680 15.680 ;
        RECT 0.000 14.840 3.640 15.120 ;
      LAYER met1 ;
        RECT 3.640 14.840 5.320 15.120 ;
      LAYER met1 ;
        RECT 5.320 14.840 6.720 15.120 ;
      LAYER met1 ;
        RECT 6.720 14.840 7.840 15.120 ;
      LAYER met1 ;
        RECT 7.840 14.840 15.680 15.120 ;
      LAYER met1 ;
        RECT 15.680 14.840 17.920 15.680 ;
      LAYER met1 ;
        RECT 17.920 15.400 30.240 15.680 ;
      LAYER met1 ;
        RECT 30.240 15.400 31.920 15.680 ;
      LAYER met1 ;
        RECT 31.920 15.400 35.840 15.680 ;
        RECT 17.920 15.120 25.480 15.400 ;
      LAYER met1 ;
        RECT 25.480 15.120 26.600 15.400 ;
      LAYER met1 ;
        RECT 26.600 15.120 30.240 15.400 ;
        RECT 17.920 14.840 24.920 15.120 ;
      LAYER met1 ;
        RECT 24.920 14.840 26.600 15.120 ;
      LAYER met1 ;
        RECT 26.600 14.840 27.440 15.120 ;
      LAYER met1 ;
        RECT 27.440 14.840 28.560 15.120 ;
      LAYER met1 ;
        RECT 0.000 14.560 3.920 14.840 ;
      LAYER met1 ;
        RECT 3.920 14.560 5.320 14.840 ;
      LAYER met1 ;
        RECT 5.320 14.560 6.440 14.840 ;
      LAYER met1 ;
        RECT 6.440 14.560 8.120 14.840 ;
      LAYER met1 ;
        RECT 8.120 14.560 24.640 14.840 ;
      LAYER met1 ;
        RECT 24.640 14.560 26.600 14.840 ;
      LAYER met1 ;
        RECT 26.600 14.560 27.160 14.840 ;
      LAYER met1 ;
        RECT 27.160 14.560 28.560 14.840 ;
      LAYER met1 ;
        RECT 28.560 14.560 30.240 15.120 ;
      LAYER met1 ;
        RECT 30.240 14.840 31.640 15.400 ;
      LAYER met1 ;
        RECT 31.640 14.840 35.840 15.400 ;
      LAYER met1 ;
        RECT 30.240 14.560 31.920 14.840 ;
      LAYER met1 ;
        RECT 31.920 14.560 35.840 14.840 ;
        RECT 0.000 14.280 4.200 14.560 ;
      LAYER met1 ;
        RECT 4.200 14.280 5.320 14.560 ;
      LAYER met1 ;
        RECT 5.320 14.280 5.880 14.560 ;
      LAYER met1 ;
        RECT 5.880 14.280 8.120 14.560 ;
      LAYER met1 ;
        RECT 8.120 14.280 9.240 14.560 ;
      LAYER met1 ;
        RECT 9.240 14.280 10.080 14.560 ;
      LAYER met1 ;
        RECT 10.080 14.280 24.360 14.560 ;
      LAYER met1 ;
        RECT 24.360 14.280 28.560 14.560 ;
      LAYER met1 ;
        RECT 28.560 14.280 30.520 14.560 ;
      LAYER met1 ;
        RECT 30.520 14.280 32.200 14.560 ;
      LAYER met1 ;
        RECT 32.200 14.280 35.840 14.560 ;
        RECT 0.000 13.720 3.920 14.280 ;
      LAYER met1 ;
        RECT 3.920 14.000 5.320 14.280 ;
      LAYER met1 ;
        RECT 5.320 14.000 5.600 14.280 ;
      LAYER met1 ;
        RECT 5.600 14.000 8.400 14.280 ;
      LAYER met1 ;
        RECT 8.400 14.000 8.960 14.280 ;
      LAYER met1 ;
        RECT 8.960 14.000 10.080 14.280 ;
        RECT 3.920 13.720 5.040 14.000 ;
      LAYER met1 ;
        RECT 0.000 13.160 3.640 13.720 ;
      LAYER met1 ;
        RECT 3.640 13.440 5.040 13.720 ;
      LAYER met1 ;
        RECT 5.040 13.440 5.600 14.000 ;
      LAYER met1 ;
        RECT 5.600 13.720 7.000 14.000 ;
      LAYER met1 ;
        RECT 7.000 13.720 7.280 14.000 ;
      LAYER met1 ;
        RECT 5.600 13.440 6.720 13.720 ;
      LAYER met1 ;
        RECT 6.720 13.440 7.280 13.720 ;
      LAYER met1 ;
        RECT 7.280 13.440 10.080 14.000 ;
      LAYER met1 ;
        RECT 10.080 13.720 24.080 14.280 ;
      LAYER met1 ;
        RECT 24.080 14.000 28.280 14.280 ;
      LAYER met1 ;
        RECT 28.280 14.000 30.800 14.280 ;
      LAYER met1 ;
        RECT 30.800 14.000 32.480 14.280 ;
        RECT 24.080 13.720 25.480 14.000 ;
      LAYER met1 ;
        RECT 25.480 13.720 25.760 14.000 ;
      LAYER met1 ;
        RECT 25.760 13.720 28.000 14.000 ;
      LAYER met1 ;
        RECT 28.000 13.720 31.080 14.000 ;
      LAYER met1 ;
        RECT 31.080 13.720 32.480 14.000 ;
      LAYER met1 ;
        RECT 32.480 13.720 35.840 14.280 ;
        RECT 10.080 13.440 20.720 13.720 ;
      LAYER met1 ;
        RECT 20.720 13.440 21.560 13.720 ;
      LAYER met1 ;
        RECT 21.560 13.440 24.080 13.720 ;
      LAYER met1 ;
        RECT 24.080 13.440 25.200 13.720 ;
      LAYER met1 ;
        RECT 25.200 13.440 25.760 13.720 ;
      LAYER met1 ;
        RECT 25.760 13.440 27.440 13.720 ;
      LAYER met1 ;
        RECT 27.440 13.440 31.360 13.720 ;
      LAYER met1 ;
        RECT 31.360 13.440 32.760 13.720 ;
      LAYER met1 ;
        RECT 32.760 13.440 35.840 13.720 ;
      LAYER met1 ;
        RECT 3.640 13.160 4.760 13.440 ;
      LAYER met1 ;
        RECT 0.000 10.640 3.360 13.160 ;
      LAYER met1 ;
        RECT 3.360 12.880 4.760 13.160 ;
      LAYER met1 ;
        RECT 4.760 12.880 7.560 13.440 ;
      LAYER met1 ;
        RECT 7.560 13.160 9.800 13.440 ;
      LAYER met1 ;
        RECT 9.800 13.160 17.080 13.440 ;
      LAYER met1 ;
        RECT 17.080 13.160 17.920 13.440 ;
      LAYER met1 ;
        RECT 17.920 13.160 20.160 13.440 ;
      LAYER met1 ;
        RECT 20.160 13.160 21.560 13.440 ;
        RECT 7.560 12.880 9.240 13.160 ;
      LAYER met1 ;
        RECT 9.240 12.880 16.800 13.160 ;
      LAYER met1 ;
        RECT 16.800 12.880 18.200 13.160 ;
      LAYER met1 ;
        RECT 18.200 12.880 19.880 13.160 ;
      LAYER met1 ;
        RECT 19.880 12.880 21.560 13.160 ;
      LAYER met1 ;
        RECT 21.560 12.880 25.760 13.440 ;
      LAYER met1 ;
        RECT 25.760 13.160 27.160 13.440 ;
      LAYER met1 ;
        RECT 27.160 13.160 31.640 13.440 ;
      LAYER met1 ;
        RECT 25.760 12.880 26.880 13.160 ;
      LAYER met1 ;
        RECT 26.880 12.880 31.640 13.160 ;
      LAYER met1 ;
        RECT 31.640 12.880 33.040 13.440 ;
      LAYER met1 ;
        RECT 33.040 12.880 35.840 13.440 ;
      LAYER met1 ;
        RECT 3.360 12.320 4.480 12.880 ;
      LAYER met1 ;
        RECT 4.480 12.600 16.520 12.880 ;
      LAYER met1 ;
        RECT 16.520 12.600 21.560 12.880 ;
      LAYER met1 ;
        RECT 21.560 12.600 31.920 12.880 ;
        RECT 4.480 12.320 14.000 12.600 ;
      LAYER met1 ;
        RECT 14.000 12.320 15.400 12.600 ;
      LAYER met1 ;
        RECT 15.400 12.320 15.960 12.600 ;
      LAYER met1 ;
        RECT 15.960 12.320 21.000 12.600 ;
      LAYER met1 ;
        RECT 21.000 12.320 31.920 12.600 ;
      LAYER met1 ;
        RECT 31.920 12.320 33.320 12.880 ;
        RECT 3.360 11.480 4.200 12.320 ;
      LAYER met1 ;
        RECT 4.200 11.760 14.000 12.320 ;
      LAYER met1 ;
        RECT 14.000 12.040 20.720 12.320 ;
      LAYER met1 ;
        RECT 20.720 12.040 31.360 12.320 ;
      LAYER met1 ;
        RECT 31.360 12.040 33.320 12.320 ;
      LAYER met1 ;
        RECT 33.320 12.040 35.840 12.880 ;
      LAYER met1 ;
        RECT 14.000 11.760 17.360 12.040 ;
      LAYER met1 ;
        RECT 17.360 11.760 18.200 12.040 ;
      LAYER met1 ;
        RECT 18.200 11.760 19.880 12.040 ;
      LAYER met1 ;
        RECT 19.880 11.760 26.880 12.040 ;
      LAYER met1 ;
        RECT 26.880 11.760 28.000 12.040 ;
      LAYER met1 ;
        RECT 28.000 11.760 30.800 12.040 ;
      LAYER met1 ;
        RECT 30.800 11.760 33.040 12.040 ;
      LAYER met1 ;
        RECT 33.040 11.760 35.840 12.040 ;
        RECT 4.200 11.480 14.560 11.760 ;
      LAYER met1 ;
        RECT 14.560 11.480 16.800 11.760 ;
      LAYER met1 ;
        RECT 16.800 11.480 26.600 11.760 ;
      LAYER met1 ;
        RECT 26.600 11.480 28.000 11.760 ;
      LAYER met1 ;
        RECT 28.000 11.480 29.120 11.760 ;
      LAYER met1 ;
        RECT 29.120 11.480 32.760 11.760 ;
      LAYER met1 ;
        RECT 32.760 11.480 35.840 11.760 ;
      LAYER met1 ;
        RECT 3.360 11.200 5.040 11.480 ;
      LAYER met1 ;
        RECT 5.040 11.200 6.440 11.480 ;
      LAYER met1 ;
        RECT 6.440 11.200 8.680 11.480 ;
      LAYER met1 ;
        RECT 8.680 11.200 26.320 11.480 ;
      LAYER met1 ;
        RECT 26.320 11.200 32.200 11.480 ;
      LAYER met1 ;
        RECT 32.200 11.200 35.840 11.480 ;
      LAYER met1 ;
        RECT 3.360 10.920 9.240 11.200 ;
      LAYER met1 ;
        RECT 9.240 10.920 25.760 11.200 ;
      LAYER met1 ;
        RECT 25.760 10.920 27.720 11.200 ;
      LAYER met1 ;
        RECT 27.720 10.920 28.000 11.200 ;
      LAYER met1 ;
        RECT 28.000 10.920 31.360 11.200 ;
      LAYER met1 ;
        RECT 31.360 10.920 35.840 11.200 ;
      LAYER met1 ;
        RECT 3.360 10.640 9.520 10.920 ;
      LAYER met1 ;
        RECT 9.520 10.640 25.200 10.920 ;
      LAYER met1 ;
        RECT 25.200 10.640 27.440 10.920 ;
      LAYER met1 ;
        RECT 27.440 10.640 28.000 10.920 ;
      LAYER met1 ;
        RECT 28.000 10.640 29.960 10.920 ;
      LAYER met1 ;
        RECT 29.960 10.640 35.840 10.920 ;
        RECT 0.000 10.360 4.200 10.640 ;
      LAYER met1 ;
        RECT 4.200 10.360 7.280 10.640 ;
      LAYER met1 ;
        RECT 7.280 10.360 7.840 10.640 ;
      LAYER met1 ;
        RECT 7.840 10.360 10.080 10.640 ;
      LAYER met1 ;
        RECT 10.080 10.360 24.640 10.640 ;
      LAYER met1 ;
        RECT 24.640 10.360 27.160 10.640 ;
      LAYER met1 ;
        RECT 27.160 10.360 35.840 10.640 ;
        RECT 0.000 10.080 8.400 10.360 ;
      LAYER met1 ;
        RECT 8.400 10.080 10.640 10.360 ;
      LAYER met1 ;
        RECT 10.640 10.080 23.800 10.360 ;
      LAYER met1 ;
        RECT 23.800 10.080 26.600 10.360 ;
      LAYER met1 ;
        RECT 26.600 10.080 35.840 10.360 ;
        RECT 0.000 9.800 8.680 10.080 ;
      LAYER met1 ;
        RECT 8.680 9.800 12.880 10.080 ;
      LAYER met1 ;
        RECT 12.880 9.800 22.960 10.080 ;
      LAYER met1 ;
        RECT 22.960 9.800 26.040 10.080 ;
      LAYER met1 ;
        RECT 26.040 9.800 35.840 10.080 ;
        RECT 0.000 9.520 9.240 9.800 ;
      LAYER met1 ;
        RECT 9.240 9.520 13.440 9.800 ;
      LAYER met1 ;
        RECT 13.440 9.520 22.960 9.800 ;
      LAYER met1 ;
        RECT 22.960 9.520 25.200 9.800 ;
      LAYER met1 ;
        RECT 25.200 9.520 35.840 9.800 ;
        RECT 0.000 9.240 9.800 9.520 ;
      LAYER met1 ;
        RECT 9.800 9.240 15.120 9.520 ;
      LAYER met1 ;
        RECT 15.120 9.240 22.960 9.520 ;
      LAYER met1 ;
        RECT 22.960 9.240 24.360 9.520 ;
      LAYER met1 ;
        RECT 24.360 9.240 35.840 9.520 ;
        RECT 0.000 8.680 10.360 9.240 ;
      LAYER met1 ;
        RECT 10.360 8.960 11.480 9.240 ;
      LAYER met1 ;
        RECT 11.480 8.960 12.040 9.240 ;
      LAYER met1 ;
        RECT 12.040 8.960 15.120 9.240 ;
      LAYER met1 ;
        RECT 15.120 8.960 35.840 9.240 ;
      LAYER met1 ;
        RECT 10.360 8.680 11.760 8.960 ;
      LAYER met1 ;
        RECT 11.760 8.680 12.880 8.960 ;
      LAYER met1 ;
        RECT 12.880 8.680 15.120 8.960 ;
      LAYER met1 ;
        RECT 15.120 8.680 24.080 8.960 ;
        RECT 0.000 8.120 10.640 8.680 ;
      LAYER met1 ;
        RECT 10.640 8.400 11.760 8.680 ;
      LAYER met1 ;
        RECT 11.760 8.400 24.080 8.680 ;
      LAYER met1 ;
        RECT 24.080 8.400 25.200 8.960 ;
      LAYER met1 ;
        RECT 25.200 8.400 35.840 8.960 ;
      LAYER met1 ;
        RECT 10.640 8.120 12.040 8.400 ;
      LAYER met1 ;
        RECT 12.040 8.120 24.080 8.400 ;
      LAYER met1 ;
        RECT 24.080 8.120 25.480 8.400 ;
      LAYER met1 ;
        RECT 25.480 8.120 35.840 8.400 ;
        RECT 0.000 7.560 10.920 8.120 ;
      LAYER met1 ;
        RECT 10.920 7.840 12.320 8.120 ;
      LAYER met1 ;
        RECT 12.320 7.840 24.360 8.120 ;
      LAYER met1 ;
        RECT 10.920 7.560 12.600 7.840 ;
      LAYER met1 ;
        RECT 12.600 7.560 24.360 7.840 ;
      LAYER met1 ;
        RECT 24.360 7.560 25.760 8.120 ;
      LAYER met1 ;
        RECT 0.000 7.280 11.200 7.560 ;
      LAYER met1 ;
        RECT 11.200 7.280 12.880 7.560 ;
      LAYER met1 ;
        RECT 12.880 7.280 24.640 7.560 ;
      LAYER met1 ;
        RECT 24.640 7.280 25.760 7.560 ;
      LAYER met1 ;
        RECT 25.760 7.280 35.840 8.120 ;
        RECT 0.000 7.000 11.480 7.280 ;
      LAYER met1 ;
        RECT 11.480 7.000 13.160 7.280 ;
      LAYER met1 ;
        RECT 0.000 6.720 11.760 7.000 ;
      LAYER met1 ;
        RECT 11.760 6.720 13.160 7.000 ;
      LAYER met1 ;
        RECT 13.160 6.720 24.920 7.280 ;
      LAYER met1 ;
        RECT 24.920 6.720 26.040 7.280 ;
      LAYER met1 ;
        RECT 26.040 6.720 35.840 7.280 ;
        RECT 0.000 6.440 12.040 6.720 ;
      LAYER met1 ;
        RECT 12.040 6.440 13.160 6.720 ;
      LAYER met1 ;
        RECT 0.000 5.880 11.760 6.440 ;
      LAYER met1 ;
        RECT 11.760 5.880 13.160 6.440 ;
      LAYER met1 ;
        RECT 13.160 5.880 25.200 6.720 ;
      LAYER met1 ;
        RECT 25.200 5.880 26.320 6.720 ;
      LAYER met1 ;
        RECT 0.000 5.600 11.480 5.880 ;
      LAYER met1 ;
        RECT 11.480 5.600 12.880 5.880 ;
      LAYER met1 ;
        RECT 12.880 5.600 25.480 5.880 ;
      LAYER met1 ;
        RECT 25.480 5.600 26.320 5.880 ;
      LAYER met1 ;
        RECT 26.320 5.600 35.840 6.720 ;
        RECT 0.000 5.320 11.200 5.600 ;
      LAYER met1 ;
        RECT 11.200 5.320 12.600 5.600 ;
      LAYER met1 ;
        RECT 12.600 5.320 25.480 5.600 ;
        RECT 0.000 5.040 10.920 5.320 ;
      LAYER met1 ;
        RECT 10.920 5.040 12.320 5.320 ;
      LAYER met1 ;
        RECT 0.000 3.920 10.640 5.040 ;
      LAYER met1 ;
        RECT 10.640 4.760 12.320 5.040 ;
      LAYER met1 ;
        RECT 12.320 4.760 25.480 5.320 ;
      LAYER met1 ;
        RECT 25.480 4.760 26.600 5.600 ;
      LAYER met1 ;
        RECT 26.600 4.760 35.840 5.600 ;
      LAYER met1 ;
        RECT 10.640 4.480 13.720 4.760 ;
      LAYER met1 ;
        RECT 13.720 4.480 25.760 4.760 ;
      LAYER met1 ;
        RECT 10.640 3.920 14.000 4.480 ;
      LAYER met1 ;
        RECT 14.000 3.920 25.760 4.480 ;
      LAYER met1 ;
        RECT 25.760 3.920 26.880 4.760 ;
      LAYER met1 ;
        RECT 0.000 3.080 12.600 3.920 ;
      LAYER met1 ;
        RECT 12.600 3.640 14.000 3.920 ;
      LAYER met1 ;
        RECT 14.000 3.640 26.040 3.920 ;
      LAYER met1 ;
        RECT 26.040 3.640 26.880 3.920 ;
      LAYER met1 ;
        RECT 26.880 3.640 35.840 4.760 ;
      LAYER met1 ;
        RECT 12.600 3.080 13.720 3.640 ;
      LAYER met1 ;
        RECT 13.720 3.080 26.040 3.640 ;
      LAYER met1 ;
        RECT 26.040 3.080 27.160 3.640 ;
      LAYER met1 ;
        RECT 0.000 2.240 12.320 3.080 ;
      LAYER met1 ;
        RECT 12.320 2.520 13.440 3.080 ;
      LAYER met1 ;
        RECT 13.440 2.520 26.320 3.080 ;
      LAYER met1 ;
        RECT 26.320 2.520 27.160 3.080 ;
      LAYER met1 ;
        RECT 27.160 2.520 35.840 3.640 ;
      LAYER met1 ;
        RECT 12.320 2.240 13.160 2.520 ;
      LAYER met1 ;
        RECT 0.000 0.280 12.040 2.240 ;
      LAYER met1 ;
        RECT 12.040 1.680 13.160 2.240 ;
      LAYER met1 ;
        RECT 13.160 1.680 26.320 2.520 ;
      LAYER met1 ;
        RECT 26.320 1.680 27.440 2.520 ;
        RECT 12.040 0.280 12.880 1.680 ;
      LAYER met1 ;
        RECT 12.880 0.280 26.600 1.680 ;
      LAYER met1 ;
        RECT 26.600 0.280 27.440 1.680 ;
      LAYER met1 ;
        RECT 27.440 0.280 35.840 2.520 ;
        RECT 0.000 0.000 35.840 0.280 ;
      LAYER met2 ;
        RECT 0.000 35.560 35.840 35.840 ;
        RECT 0.000 35.280 29.960 35.560 ;
      LAYER met2 ;
        RECT 29.960 35.280 31.360 35.560 ;
      LAYER met2 ;
        RECT 0.000 34.160 4.200 35.280 ;
      LAYER met2 ;
        RECT 4.200 35.000 5.600 35.280 ;
      LAYER met2 ;
        RECT 5.600 35.000 29.120 35.280 ;
      LAYER met2 ;
        RECT 29.120 35.000 31.360 35.280 ;
      LAYER met2 ;
        RECT 31.360 35.000 35.840 35.560 ;
      LAYER met2 ;
        RECT 4.200 34.720 6.720 35.000 ;
      LAYER met2 ;
        RECT 6.720 34.720 28.560 35.000 ;
      LAYER met2 ;
        RECT 28.560 34.720 31.640 35.000 ;
        RECT 4.200 34.440 7.560 34.720 ;
      LAYER met2 ;
        RECT 7.560 34.440 27.720 34.720 ;
      LAYER met2 ;
        RECT 27.720 34.440 31.640 34.720 ;
        RECT 4.200 34.160 8.120 34.440 ;
      LAYER met2 ;
        RECT 8.120 34.160 27.160 34.440 ;
      LAYER met2 ;
        RECT 27.160 34.160 29.960 34.440 ;
      LAYER met2 ;
        RECT 29.960 34.160 30.800 34.440 ;
      LAYER met2 ;
        RECT 30.800 34.160 31.640 34.440 ;
      LAYER met2 ;
        RECT 31.640 34.160 35.840 35.000 ;
        RECT 0.000 33.040 3.920 34.160 ;
      LAYER met2 ;
        RECT 3.920 33.320 5.040 34.160 ;
      LAYER met2 ;
        RECT 5.040 33.880 6.160 34.160 ;
      LAYER met2 ;
        RECT 6.160 33.880 8.400 34.160 ;
      LAYER met2 ;
        RECT 8.400 33.880 26.600 34.160 ;
      LAYER met2 ;
        RECT 26.600 33.880 29.120 34.160 ;
      LAYER met2 ;
        RECT 29.120 33.880 30.800 34.160 ;
        RECT 5.040 33.600 6.720 33.880 ;
      LAYER met2 ;
        RECT 6.720 33.600 8.680 33.880 ;
      LAYER met2 ;
        RECT 8.680 33.600 26.040 33.880 ;
      LAYER met2 ;
        RECT 26.040 33.600 28.560 33.880 ;
      LAYER met2 ;
        RECT 28.560 33.600 30.800 33.880 ;
      LAYER met2 ;
        RECT 30.800 33.600 31.920 34.160 ;
      LAYER met2 ;
        RECT 5.040 33.320 7.280 33.600 ;
      LAYER met2 ;
        RECT 7.280 33.320 8.960 33.600 ;
      LAYER met2 ;
        RECT 8.960 33.320 25.760 33.600 ;
      LAYER met2 ;
        RECT 25.760 33.320 28.000 33.600 ;
      LAYER met2 ;
        RECT 28.000 33.320 31.080 33.600 ;
      LAYER met2 ;
        RECT 31.080 33.320 31.920 33.600 ;
      LAYER met2 ;
        RECT 31.920 33.320 35.840 34.160 ;
      LAYER met2 ;
        RECT 3.920 33.040 4.760 33.320 ;
      LAYER met2 ;
        RECT 4.760 33.040 7.560 33.320 ;
      LAYER met2 ;
        RECT 7.560 33.040 9.240 33.320 ;
      LAYER met2 ;
        RECT 9.240 33.040 13.720 33.320 ;
      LAYER met2 ;
        RECT 13.720 33.040 14.560 33.320 ;
      LAYER met2 ;
        RECT 14.560 33.040 25.200 33.320 ;
      LAYER met2 ;
        RECT 25.200 33.040 27.440 33.320 ;
      LAYER met2 ;
        RECT 27.440 33.040 31.080 33.320 ;
        RECT 0.000 31.640 3.640 33.040 ;
      LAYER met2 ;
        RECT 3.640 32.480 4.760 33.040 ;
      LAYER met2 ;
        RECT 4.760 32.760 7.840 33.040 ;
      LAYER met2 ;
        RECT 7.840 32.760 9.800 33.040 ;
      LAYER met2 ;
        RECT 9.800 32.760 13.720 33.040 ;
      LAYER met2 ;
        RECT 13.720 32.760 16.800 33.040 ;
      LAYER met2 ;
        RECT 16.800 32.760 24.920 33.040 ;
      LAYER met2 ;
        RECT 24.920 32.760 26.880 33.040 ;
      LAYER met2 ;
        RECT 26.880 32.760 31.080 33.040 ;
      LAYER met2 ;
        RECT 31.080 32.760 32.200 33.320 ;
      LAYER met2 ;
        RECT 4.760 32.480 8.400 32.760 ;
      LAYER met2 ;
        RECT 8.400 32.480 10.080 32.760 ;
      LAYER met2 ;
        RECT 10.080 32.480 13.720 32.760 ;
      LAYER met2 ;
        RECT 13.720 32.480 17.640 32.760 ;
      LAYER met2 ;
        RECT 17.640 32.480 24.640 32.760 ;
      LAYER met2 ;
        RECT 24.640 32.480 26.320 32.760 ;
      LAYER met2 ;
        RECT 26.320 32.480 31.360 32.760 ;
      LAYER met2 ;
        RECT 31.360 32.480 32.200 32.760 ;
      LAYER met2 ;
        RECT 32.200 32.480 35.840 33.320 ;
      LAYER met2 ;
        RECT 3.640 31.640 4.480 32.480 ;
      LAYER met2 ;
        RECT 4.480 32.200 8.680 32.480 ;
      LAYER met2 ;
        RECT 8.680 32.200 10.640 32.480 ;
      LAYER met2 ;
        RECT 10.640 32.200 13.720 32.480 ;
      LAYER met2 ;
        RECT 13.720 32.200 18.480 32.480 ;
      LAYER met2 ;
        RECT 18.480 32.200 24.080 32.480 ;
      LAYER met2 ;
        RECT 24.080 32.200 26.040 32.480 ;
      LAYER met2 ;
        RECT 26.040 32.200 31.360 32.480 ;
        RECT 4.480 31.920 8.960 32.200 ;
      LAYER met2 ;
        RECT 8.960 31.920 10.920 32.200 ;
      LAYER met2 ;
        RECT 10.920 31.920 13.720 32.200 ;
      LAYER met2 ;
        RECT 13.720 31.920 14.840 32.200 ;
      LAYER met2 ;
        RECT 14.840 31.920 15.960 32.200 ;
      LAYER met2 ;
        RECT 15.960 31.920 19.320 32.200 ;
      LAYER met2 ;
        RECT 19.320 31.920 23.800 32.200 ;
      LAYER met2 ;
        RECT 23.800 31.920 25.760 32.200 ;
      LAYER met2 ;
        RECT 25.760 31.920 31.360 32.200 ;
        RECT 4.480 31.640 9.520 31.920 ;
      LAYER met2 ;
        RECT 9.520 31.640 11.200 31.920 ;
      LAYER met2 ;
        RECT 11.200 31.640 14.000 31.920 ;
      LAYER met2 ;
        RECT 14.000 31.640 14.840 31.920 ;
      LAYER met2 ;
        RECT 14.840 31.640 17.080 31.920 ;
      LAYER met2 ;
        RECT 17.080 31.640 19.880 31.920 ;
      LAYER met2 ;
        RECT 19.880 31.640 23.800 31.920 ;
      LAYER met2 ;
        RECT 23.800 31.640 25.480 31.920 ;
      LAYER met2 ;
        RECT 25.480 31.640 31.360 31.920 ;
      LAYER met2 ;
        RECT 31.360 31.640 32.480 32.480 ;
      LAYER met2 ;
        RECT 0.000 30.240 3.360 31.640 ;
      LAYER met2 ;
        RECT 3.360 31.080 4.480 31.640 ;
      LAYER met2 ;
        RECT 4.480 31.360 9.800 31.640 ;
      LAYER met2 ;
        RECT 9.800 31.360 11.480 31.640 ;
      LAYER met2 ;
        RECT 11.480 31.360 14.000 31.640 ;
        RECT 4.480 31.080 10.080 31.360 ;
      LAYER met2 ;
        RECT 10.080 31.080 11.760 31.360 ;
      LAYER met2 ;
        RECT 11.760 31.080 14.000 31.360 ;
      LAYER met2 ;
        RECT 14.000 31.080 15.120 31.640 ;
      LAYER met2 ;
        RECT 15.120 31.360 17.920 31.640 ;
      LAYER met2 ;
        RECT 17.920 31.360 20.440 31.640 ;
      LAYER met2 ;
        RECT 20.440 31.360 23.520 31.640 ;
      LAYER met2 ;
        RECT 23.520 31.360 25.200 31.640 ;
      LAYER met2 ;
        RECT 25.200 31.360 31.640 31.640 ;
      LAYER met2 ;
        RECT 31.640 31.360 32.480 31.640 ;
      LAYER met2 ;
        RECT 32.480 31.360 35.840 32.480 ;
        RECT 15.120 31.080 18.480 31.360 ;
      LAYER met2 ;
        RECT 18.480 31.080 21.000 31.360 ;
      LAYER met2 ;
        RECT 21.000 31.080 23.520 31.360 ;
      LAYER met2 ;
        RECT 23.520 31.080 24.920 31.360 ;
      LAYER met2 ;
        RECT 24.920 31.080 31.640 31.360 ;
      LAYER met2 ;
        RECT 3.360 30.240 4.200 31.080 ;
      LAYER met2 ;
        RECT 4.200 30.800 10.360 31.080 ;
      LAYER met2 ;
        RECT 10.360 30.800 12.040 31.080 ;
      LAYER met2 ;
        RECT 4.200 30.520 10.640 30.800 ;
      LAYER met2 ;
        RECT 10.640 30.520 12.040 30.800 ;
      LAYER met2 ;
        RECT 12.040 30.520 14.280 31.080 ;
      LAYER met2 ;
        RECT 14.280 30.520 15.400 31.080 ;
      LAYER met2 ;
        RECT 15.400 30.800 19.040 31.080 ;
      LAYER met2 ;
        RECT 19.040 30.800 21.280 31.080 ;
      LAYER met2 ;
        RECT 21.280 30.800 23.240 31.080 ;
      LAYER met2 ;
        RECT 23.240 30.800 24.360 31.080 ;
      LAYER met2 ;
        RECT 15.400 30.520 19.600 30.800 ;
      LAYER met2 ;
        RECT 19.600 30.520 21.560 30.800 ;
      LAYER met2 ;
        RECT 21.560 30.520 22.960 30.800 ;
      LAYER met2 ;
        RECT 22.960 30.520 24.360 30.800 ;
      LAYER met2 ;
        RECT 24.360 30.520 31.640 31.080 ;
      LAYER met2 ;
        RECT 31.640 30.520 32.760 31.360 ;
      LAYER met2 ;
        RECT 4.200 30.240 10.920 30.520 ;
      LAYER met2 ;
        RECT 10.920 30.240 12.320 30.520 ;
      LAYER met2 ;
        RECT 12.320 30.240 14.280 30.520 ;
      LAYER met2 ;
        RECT 14.280 30.240 15.680 30.520 ;
      LAYER met2 ;
        RECT 15.680 30.240 20.160 30.520 ;
      LAYER met2 ;
        RECT 20.160 30.240 21.840 30.520 ;
      LAYER met2 ;
        RECT 21.840 30.240 22.960 30.520 ;
      LAYER met2 ;
        RECT 22.960 30.240 24.080 30.520 ;
      LAYER met2 ;
        RECT 0.000 28.000 3.080 30.240 ;
      LAYER met2 ;
        RECT 3.080 29.680 4.200 30.240 ;
      LAYER met2 ;
        RECT 4.200 29.960 11.200 30.240 ;
      LAYER met2 ;
        RECT 11.200 29.960 12.600 30.240 ;
      LAYER met2 ;
        RECT 12.600 29.960 14.560 30.240 ;
      LAYER met2 ;
        RECT 14.560 29.960 15.960 30.240 ;
      LAYER met2 ;
        RECT 15.960 29.960 20.440 30.240 ;
      LAYER met2 ;
        RECT 20.440 29.960 22.400 30.240 ;
      LAYER met2 ;
        RECT 22.400 29.960 22.680 30.240 ;
      LAYER met2 ;
        RECT 22.680 29.960 24.080 30.240 ;
      LAYER met2 ;
        RECT 24.080 29.960 31.920 30.520 ;
      LAYER met2 ;
        RECT 31.920 29.960 32.760 30.520 ;
      LAYER met2 ;
        RECT 32.760 29.960 35.840 31.360 ;
        RECT 4.200 29.680 11.480 29.960 ;
      LAYER met2 ;
        RECT 11.480 29.680 12.880 29.960 ;
      LAYER met2 ;
        RECT 12.880 29.680 14.560 29.960 ;
      LAYER met2 ;
        RECT 14.560 29.680 16.240 29.960 ;
      LAYER met2 ;
        RECT 16.240 29.680 21.000 29.960 ;
      LAYER met2 ;
        RECT 21.000 29.680 23.800 29.960 ;
        RECT 3.080 28.000 3.920 29.680 ;
      LAYER met2 ;
        RECT 3.920 29.400 11.760 29.680 ;
      LAYER met2 ;
        RECT 11.760 29.400 13.160 29.680 ;
      LAYER met2 ;
        RECT 13.160 29.400 14.840 29.680 ;
      LAYER met2 ;
        RECT 14.840 29.400 16.520 29.680 ;
      LAYER met2 ;
        RECT 16.520 29.400 21.280 29.680 ;
      LAYER met2 ;
        RECT 21.280 29.400 23.800 29.680 ;
      LAYER met2 ;
        RECT 23.800 29.400 31.920 29.960 ;
      LAYER met2 ;
        RECT 31.920 29.400 33.040 29.960 ;
      LAYER met2 ;
        RECT 3.920 29.120 12.040 29.400 ;
      LAYER met2 ;
        RECT 12.040 29.120 13.440 29.400 ;
      LAYER met2 ;
        RECT 13.440 29.120 15.120 29.400 ;
      LAYER met2 ;
        RECT 15.120 29.120 16.520 29.400 ;
      LAYER met2 ;
        RECT 16.520 29.120 21.560 29.400 ;
      LAYER met2 ;
        RECT 21.560 29.120 23.520 29.400 ;
      LAYER met2 ;
        RECT 3.920 28.560 12.320 29.120 ;
      LAYER met2 ;
        RECT 12.320 28.840 13.720 29.120 ;
      LAYER met2 ;
        RECT 13.720 28.840 15.400 29.120 ;
      LAYER met2 ;
        RECT 15.400 28.840 16.800 29.120 ;
      LAYER met2 ;
        RECT 16.800 28.840 21.840 29.120 ;
      LAYER met2 ;
        RECT 21.840 28.840 23.520 29.120 ;
      LAYER met2 ;
        RECT 23.520 28.840 32.200 29.400 ;
      LAYER met2 ;
        RECT 32.200 28.840 33.040 29.400 ;
      LAYER met2 ;
        RECT 33.040 28.840 35.840 29.960 ;
      LAYER met2 ;
        RECT 12.320 28.560 14.000 28.840 ;
      LAYER met2 ;
        RECT 14.000 28.560 14.560 28.840 ;
      LAYER met2 ;
        RECT 14.560 28.560 16.800 28.840 ;
      LAYER met2 ;
        RECT 16.800 28.560 22.120 28.840 ;
      LAYER met2 ;
        RECT 22.120 28.560 23.240 28.840 ;
      LAYER met2 ;
        RECT 3.920 28.280 12.600 28.560 ;
      LAYER met2 ;
        RECT 12.600 28.280 16.800 28.560 ;
      LAYER met2 ;
        RECT 16.800 28.280 22.400 28.560 ;
        RECT 3.920 28.000 12.880 28.280 ;
      LAYER met2 ;
        RECT 12.880 28.000 16.240 28.280 ;
      LAYER met2 ;
        RECT 16.240 28.000 22.400 28.280 ;
      LAYER met2 ;
        RECT 22.400 28.000 23.240 28.560 ;
      LAYER met2 ;
        RECT 23.240 28.000 32.200 28.840 ;
      LAYER met2 ;
        RECT 32.200 28.000 33.320 28.840 ;
      LAYER met2 ;
        RECT 0.000 26.320 2.800 28.000 ;
      LAYER met2 ;
        RECT 2.800 27.440 3.920 28.000 ;
      LAYER met2 ;
        RECT 3.920 27.720 13.440 28.000 ;
      LAYER met2 ;
        RECT 13.440 27.720 15.120 28.000 ;
      LAYER met2 ;
        RECT 15.120 27.720 32.480 28.000 ;
        RECT 3.920 27.440 13.160 27.720 ;
      LAYER met2 ;
        RECT 13.160 27.440 14.840 27.720 ;
      LAYER met2 ;
        RECT 14.840 27.440 32.480 27.720 ;
      LAYER met2 ;
        RECT 2.800 26.320 3.640 27.440 ;
      LAYER met2 ;
        RECT 3.640 27.160 12.880 27.440 ;
      LAYER met2 ;
        RECT 12.880 27.160 14.560 27.440 ;
      LAYER met2 ;
        RECT 14.560 27.160 32.480 27.440 ;
      LAYER met2 ;
        RECT 32.480 27.160 33.320 28.000 ;
      LAYER met2 ;
        RECT 33.320 27.160 35.840 28.840 ;
        RECT 0.000 23.800 2.520 26.320 ;
      LAYER met2 ;
        RECT 2.520 25.480 3.640 26.320 ;
      LAYER met2 ;
        RECT 3.640 26.040 12.600 27.160 ;
      LAYER met2 ;
        RECT 12.600 26.880 14.280 27.160 ;
      LAYER met2 ;
        RECT 14.280 26.880 32.480 27.160 ;
      LAYER met2 ;
        RECT 12.600 26.600 17.360 26.880 ;
      LAYER met2 ;
        RECT 17.360 26.600 32.480 26.880 ;
      LAYER met2 ;
        RECT 32.480 26.600 33.600 27.160 ;
        RECT 12.600 26.040 18.200 26.600 ;
      LAYER met2 ;
        RECT 3.640 25.760 16.520 26.040 ;
      LAYER met2 ;
        RECT 16.520 25.760 18.200 26.040 ;
      LAYER met2 ;
        RECT 18.200 25.760 32.760 26.600 ;
      LAYER met2 ;
        RECT 32.760 26.320 33.600 26.600 ;
      LAYER met2 ;
        RECT 33.600 26.320 35.840 27.160 ;
        RECT 3.640 25.480 32.760 25.760 ;
      LAYER met2 ;
        RECT 32.760 25.480 33.880 26.320 ;
      LAYER met2 ;
        RECT 33.880 25.480 35.840 26.320 ;
      LAYER met2 ;
        RECT 2.520 24.640 3.360 25.480 ;
      LAYER met2 ;
        RECT 3.360 24.640 32.760 25.480 ;
      LAYER met2 ;
        RECT 2.520 23.800 3.640 24.640 ;
      LAYER met2 ;
        RECT 3.640 24.360 32.760 24.640 ;
      LAYER met2 ;
        RECT 32.760 24.360 33.600 25.480 ;
      LAYER met2 ;
        RECT 0.000 22.680 2.800 23.800 ;
      LAYER met2 ;
        RECT 2.800 23.520 3.640 23.800 ;
      LAYER met2 ;
        RECT 3.640 23.520 32.480 24.360 ;
      LAYER met2 ;
        RECT 32.480 23.520 33.600 24.360 ;
      LAYER met2 ;
        RECT 33.600 23.520 35.840 25.480 ;
      LAYER met2 ;
        RECT 2.800 22.680 3.920 23.520 ;
      LAYER met2 ;
        RECT 3.920 22.960 32.480 23.520 ;
      LAYER met2 ;
        RECT 32.480 22.960 33.320 23.520 ;
      LAYER met2 ;
        RECT 3.920 22.680 32.200 22.960 ;
        RECT 0.000 21.840 3.080 22.680 ;
      LAYER met2 ;
        RECT 3.080 22.120 4.200 22.680 ;
      LAYER met2 ;
        RECT 4.200 22.400 32.200 22.680 ;
      LAYER met2 ;
        RECT 32.200 22.400 33.320 22.960 ;
      LAYER met2 ;
        RECT 33.320 22.400 35.840 23.520 ;
        RECT 4.200 22.120 31.920 22.400 ;
      LAYER met2 ;
        RECT 31.920 22.120 33.040 22.400 ;
        RECT 3.080 21.840 4.480 22.120 ;
      LAYER met2 ;
        RECT 4.480 21.840 31.640 22.120 ;
      LAYER met2 ;
        RECT 31.640 21.840 33.040 22.120 ;
      LAYER met2 ;
        RECT 33.040 21.840 35.840 22.400 ;
        RECT 0.000 21.280 3.360 21.840 ;
      LAYER met2 ;
        RECT 3.360 21.280 4.480 21.840 ;
      LAYER met2 ;
        RECT 4.480 21.560 22.120 21.840 ;
      LAYER met2 ;
        RECT 22.120 21.560 28.000 21.840 ;
      LAYER met2 ;
        RECT 28.000 21.560 31.640 21.840 ;
      LAYER met2 ;
        RECT 31.640 21.560 32.760 21.840 ;
      LAYER met2 ;
        RECT 4.480 21.280 21.560 21.560 ;
      LAYER met2 ;
        RECT 21.560 21.280 28.000 21.560 ;
      LAYER met2 ;
        RECT 28.000 21.280 31.360 21.560 ;
      LAYER met2 ;
        RECT 31.360 21.280 32.760 21.560 ;
      LAYER met2 ;
        RECT 32.760 21.280 35.840 21.840 ;
        RECT 0.000 20.440 3.640 21.280 ;
      LAYER met2 ;
        RECT 3.640 20.440 4.760 21.280 ;
      LAYER met2 ;
        RECT 4.760 20.440 7.560 21.280 ;
      LAYER met2 ;
        RECT 7.560 21.000 14.280 21.280 ;
      LAYER met2 ;
        RECT 14.280 21.000 21.000 21.280 ;
      LAYER met2 ;
        RECT 21.000 21.000 28.000 21.280 ;
      LAYER met2 ;
        RECT 28.000 21.000 31.080 21.280 ;
      LAYER met2 ;
        RECT 31.080 21.000 32.480 21.280 ;
        RECT 7.560 20.440 14.840 21.000 ;
      LAYER met2 ;
        RECT 14.840 20.440 21.000 21.000 ;
      LAYER met2 ;
        RECT 21.000 20.440 24.360 21.000 ;
      LAYER met2 ;
        RECT 24.360 20.440 25.760 21.000 ;
      LAYER met2 ;
        RECT 25.760 20.440 27.160 21.000 ;
      LAYER met2 ;
        RECT 27.160 20.720 30.800 21.000 ;
      LAYER met2 ;
        RECT 30.800 20.720 32.480 21.000 ;
      LAYER met2 ;
        RECT 32.480 20.720 35.840 21.280 ;
        RECT 27.160 20.440 30.520 20.720 ;
      LAYER met2 ;
        RECT 30.520 20.440 32.200 20.720 ;
      LAYER met2 ;
        RECT 32.200 20.440 35.840 20.720 ;
        RECT 0.000 19.880 3.920 20.440 ;
      LAYER met2 ;
        RECT 3.920 19.880 5.040 20.440 ;
      LAYER met2 ;
        RECT 5.040 20.160 8.400 20.440 ;
      LAYER met2 ;
        RECT 8.400 20.160 9.800 20.440 ;
      LAYER met2 ;
        RECT 5.040 19.880 8.120 20.160 ;
      LAYER met2 ;
        RECT 8.120 19.880 9.800 20.160 ;
      LAYER met2 ;
        RECT 9.800 19.880 11.200 20.440 ;
        RECT 0.000 19.040 4.200 19.880 ;
      LAYER met2 ;
        RECT 4.200 19.320 5.320 19.880 ;
      LAYER met2 ;
        RECT 5.320 19.600 8.120 19.880 ;
      LAYER met2 ;
        RECT 8.120 19.600 9.520 19.880 ;
      LAYER met2 ;
        RECT 9.520 19.600 11.200 19.880 ;
        RECT 5.320 19.320 7.840 19.600 ;
      LAYER met2 ;
        RECT 7.840 19.320 9.240 19.600 ;
      LAYER met2 ;
        RECT 9.240 19.320 11.200 19.600 ;
      LAYER met2 ;
        RECT 4.200 19.040 5.600 19.320 ;
      LAYER met2 ;
        RECT 0.000 18.760 4.480 19.040 ;
      LAYER met2 ;
        RECT 4.480 18.760 5.600 19.040 ;
      LAYER met2 ;
        RECT 5.600 18.760 7.840 19.320 ;
      LAYER met2 ;
        RECT 7.840 18.760 8.960 19.320 ;
      LAYER met2 ;
        RECT 8.960 18.760 11.200 19.320 ;
        RECT 0.000 17.360 1.680 18.760 ;
      LAYER met2 ;
        RECT 1.680 18.480 2.520 18.760 ;
      LAYER met2 ;
        RECT 2.520 18.480 4.480 18.760 ;
      LAYER met2 ;
        RECT 4.480 18.480 5.880 18.760 ;
        RECT 1.680 18.200 3.360 18.480 ;
      LAYER met2 ;
        RECT 3.360 18.200 4.760 18.480 ;
      LAYER met2 ;
        RECT 4.760 18.200 5.880 18.480 ;
      LAYER met2 ;
        RECT 5.880 18.200 7.560 18.760 ;
      LAYER met2 ;
        RECT 1.680 17.360 7.000 18.200 ;
      LAYER met2 ;
        RECT 7.000 17.360 7.560 18.200 ;
      LAYER met2 ;
        RECT 7.560 17.920 8.680 18.760 ;
      LAYER met2 ;
        RECT 8.680 17.920 11.200 18.760 ;
      LAYER met2 ;
        RECT 11.200 17.920 15.120 20.440 ;
      LAYER met2 ;
        RECT 15.120 17.920 20.720 20.440 ;
        RECT 0.000 16.800 1.960 17.360 ;
      LAYER met2 ;
        RECT 1.960 17.080 3.080 17.360 ;
      LAYER met2 ;
        RECT 3.080 17.080 7.560 17.360 ;
      LAYER met2 ;
        RECT 7.560 17.080 8.400 17.920 ;
      LAYER met2 ;
        RECT 8.400 17.080 11.200 17.920 ;
      LAYER met2 ;
        RECT 11.200 17.080 14.840 17.920 ;
      LAYER met2 ;
        RECT 14.840 17.080 20.720 17.920 ;
      LAYER met2 ;
        RECT 20.720 17.080 24.360 20.440 ;
      LAYER met2 ;
        RECT 24.360 20.160 26.040 20.440 ;
      LAYER met2 ;
        RECT 26.040 20.160 27.160 20.440 ;
      LAYER met2 ;
        RECT 27.160 20.160 30.240 20.440 ;
      LAYER met2 ;
        RECT 30.240 20.160 31.920 20.440 ;
      LAYER met2 ;
        RECT 31.920 20.160 35.840 20.440 ;
        RECT 24.360 19.600 26.320 20.160 ;
      LAYER met2 ;
        RECT 26.320 19.600 27.440 20.160 ;
      LAYER met2 ;
        RECT 27.440 19.880 30.240 20.160 ;
      LAYER met2 ;
        RECT 30.240 19.880 31.640 20.160 ;
      LAYER met2 ;
        RECT 31.640 19.880 35.840 20.160 ;
        RECT 27.440 19.600 29.680 19.880 ;
      LAYER met2 ;
        RECT 29.680 19.600 31.360 19.880 ;
      LAYER met2 ;
        RECT 31.360 19.600 35.840 19.880 ;
        RECT 24.360 18.200 26.600 19.600 ;
      LAYER met2 ;
        RECT 26.600 19.040 27.440 19.600 ;
      LAYER met2 ;
        RECT 27.440 19.320 29.400 19.600 ;
      LAYER met2 ;
        RECT 29.400 19.320 34.440 19.600 ;
      LAYER met2 ;
        RECT 27.440 19.040 29.120 19.320 ;
      LAYER met2 ;
        RECT 26.600 18.200 27.720 19.040 ;
      LAYER met2 ;
        RECT 27.720 18.200 29.120 19.040 ;
      LAYER met2 ;
        RECT 29.120 18.760 34.440 19.320 ;
        RECT 29.120 18.480 31.920 18.760 ;
      LAYER met2 ;
        RECT 31.920 18.480 33.040 18.760 ;
      LAYER met2 ;
        RECT 33.040 18.480 34.440 18.760 ;
      LAYER met2 ;
        RECT 34.440 18.480 35.840 19.600 ;
      LAYER met2 ;
        RECT 29.120 18.200 29.960 18.480 ;
      LAYER met2 ;
        RECT 29.960 18.200 32.760 18.480 ;
      LAYER met2 ;
        RECT 32.760 18.200 34.160 18.480 ;
      LAYER met2 ;
        RECT 34.160 18.200 35.840 18.480 ;
        RECT 24.360 17.360 26.880 18.200 ;
      LAYER met2 ;
        RECT 26.880 17.360 27.720 18.200 ;
      LAYER met2 ;
        RECT 27.720 17.920 32.760 18.200 ;
      LAYER met2 ;
        RECT 32.760 17.920 33.880 18.200 ;
      LAYER met2 ;
        RECT 27.720 17.640 32.480 17.920 ;
      LAYER met2 ;
        RECT 32.480 17.640 33.880 17.920 ;
      LAYER met2 ;
        RECT 33.880 17.640 35.840 18.200 ;
        RECT 27.720 17.360 32.200 17.640 ;
      LAYER met2 ;
        RECT 32.200 17.360 33.600 17.640 ;
      LAYER met2 ;
        RECT 33.600 17.360 35.840 17.640 ;
        RECT 24.360 17.080 26.600 17.360 ;
      LAYER met2 ;
        RECT 1.960 16.800 3.360 17.080 ;
      LAYER met2 ;
        RECT 3.360 16.800 7.560 17.080 ;
        RECT 0.000 16.520 2.240 16.800 ;
      LAYER met2 ;
        RECT 2.240 16.520 3.640 16.800 ;
      LAYER met2 ;
        RECT 3.640 16.520 7.560 16.800 ;
        RECT 0.000 15.960 2.520 16.520 ;
      LAYER met2 ;
        RECT 2.520 16.240 3.920 16.520 ;
      LAYER met2 ;
        RECT 3.920 16.240 7.560 16.520 ;
      LAYER met2 ;
        RECT 7.560 16.240 8.680 17.080 ;
      LAYER met2 ;
        RECT 8.680 16.520 11.480 17.080 ;
      LAYER met2 ;
        RECT 11.480 16.520 14.560 17.080 ;
      LAYER met2 ;
        RECT 14.560 16.520 21.000 17.080 ;
      LAYER met2 ;
        RECT 21.000 16.520 24.080 17.080 ;
      LAYER met2 ;
        RECT 24.080 16.520 26.600 17.080 ;
      LAYER met2 ;
        RECT 26.600 16.520 27.720 17.360 ;
      LAYER met2 ;
        RECT 27.720 17.080 31.920 17.360 ;
      LAYER met2 ;
        RECT 31.920 17.080 33.320 17.360 ;
      LAYER met2 ;
        RECT 33.320 17.080 35.840 17.360 ;
        RECT 27.720 16.800 31.640 17.080 ;
      LAYER met2 ;
        RECT 31.640 16.800 33.040 17.080 ;
      LAYER met2 ;
        RECT 33.040 16.800 35.840 17.080 ;
        RECT 27.720 16.520 31.360 16.800 ;
      LAYER met2 ;
        RECT 31.360 16.520 32.760 16.800 ;
      LAYER met2 ;
        RECT 8.680 16.240 11.760 16.520 ;
      LAYER met2 ;
        RECT 11.760 16.240 14.280 16.520 ;
      LAYER met2 ;
        RECT 14.280 16.240 21.280 16.520 ;
      LAYER met2 ;
        RECT 21.280 16.240 23.800 16.520 ;
      LAYER met2 ;
        RECT 23.800 16.240 26.600 16.520 ;
      LAYER met2 ;
        RECT 2.520 15.960 4.200 16.240 ;
      LAYER met2 ;
        RECT 4.200 15.960 7.840 16.240 ;
        RECT 0.000 15.680 2.800 15.960 ;
      LAYER met2 ;
        RECT 2.800 15.680 4.480 15.960 ;
      LAYER met2 ;
        RECT 4.480 15.680 7.840 15.960 ;
        RECT 0.000 15.400 3.080 15.680 ;
      LAYER met2 ;
        RECT 3.080 15.400 4.760 15.680 ;
      LAYER met2 ;
        RECT 4.760 15.400 7.840 15.680 ;
      LAYER met2 ;
        RECT 7.840 15.400 8.960 16.240 ;
      LAYER met2 ;
        RECT 8.960 15.960 11.760 16.240 ;
      LAYER met2 ;
        RECT 11.760 15.960 14.000 16.240 ;
      LAYER met2 ;
        RECT 14.000 15.960 21.840 16.240 ;
      LAYER met2 ;
        RECT 21.840 15.960 23.240 16.240 ;
      LAYER met2 ;
        RECT 23.240 15.960 26.600 16.240 ;
      LAYER met2 ;
        RECT 26.600 15.960 27.440 16.520 ;
      LAYER met2 ;
        RECT 27.440 16.240 31.080 16.520 ;
      LAYER met2 ;
        RECT 31.080 16.240 32.760 16.520 ;
      LAYER met2 ;
        RECT 32.760 16.240 35.840 16.800 ;
        RECT 27.440 15.960 30.800 16.240 ;
      LAYER met2 ;
        RECT 30.800 15.960 32.480 16.240 ;
      LAYER met2 ;
        RECT 32.480 15.960 35.840 16.240 ;
        RECT 8.960 15.680 12.040 15.960 ;
      LAYER met2 ;
        RECT 12.040 15.680 13.720 15.960 ;
      LAYER met2 ;
        RECT 13.720 15.680 30.520 15.960 ;
      LAYER met2 ;
        RECT 30.520 15.680 32.200 15.960 ;
      LAYER met2 ;
        RECT 32.200 15.680 35.840 15.960 ;
        RECT 0.000 15.120 3.360 15.400 ;
      LAYER met2 ;
        RECT 3.360 15.120 5.040 15.400 ;
      LAYER met2 ;
        RECT 5.040 15.120 8.120 15.400 ;
      LAYER met2 ;
        RECT 8.120 15.120 8.960 15.400 ;
      LAYER met2 ;
        RECT 8.960 15.120 15.680 15.680 ;
        RECT 0.000 14.840 3.640 15.120 ;
      LAYER met2 ;
        RECT 3.640 14.840 5.320 15.120 ;
      LAYER met2 ;
        RECT 5.320 14.840 6.720 15.120 ;
      LAYER met2 ;
        RECT 6.720 14.840 7.840 15.120 ;
      LAYER met2 ;
        RECT 7.840 14.840 15.680 15.120 ;
      LAYER met2 ;
        RECT 15.680 14.840 17.920 15.680 ;
      LAYER met2 ;
        RECT 17.920 15.400 30.240 15.680 ;
      LAYER met2 ;
        RECT 30.240 15.400 31.920 15.680 ;
      LAYER met2 ;
        RECT 31.920 15.400 35.840 15.680 ;
        RECT 17.920 15.120 25.480 15.400 ;
      LAYER met2 ;
        RECT 25.480 15.120 26.600 15.400 ;
      LAYER met2 ;
        RECT 26.600 15.120 30.240 15.400 ;
        RECT 17.920 14.840 24.920 15.120 ;
      LAYER met2 ;
        RECT 24.920 14.840 26.600 15.120 ;
      LAYER met2 ;
        RECT 26.600 14.840 27.440 15.120 ;
      LAYER met2 ;
        RECT 27.440 14.840 28.560 15.120 ;
      LAYER met2 ;
        RECT 0.000 14.560 3.920 14.840 ;
      LAYER met2 ;
        RECT 3.920 14.560 5.320 14.840 ;
      LAYER met2 ;
        RECT 5.320 14.560 6.440 14.840 ;
      LAYER met2 ;
        RECT 6.440 14.560 8.120 14.840 ;
      LAYER met2 ;
        RECT 8.120 14.560 24.640 14.840 ;
      LAYER met2 ;
        RECT 24.640 14.560 26.600 14.840 ;
      LAYER met2 ;
        RECT 26.600 14.560 27.160 14.840 ;
      LAYER met2 ;
        RECT 27.160 14.560 28.560 14.840 ;
      LAYER met2 ;
        RECT 28.560 14.560 30.240 15.120 ;
      LAYER met2 ;
        RECT 30.240 14.840 31.640 15.400 ;
      LAYER met2 ;
        RECT 31.640 14.840 35.840 15.400 ;
      LAYER met2 ;
        RECT 30.240 14.560 31.920 14.840 ;
      LAYER met2 ;
        RECT 31.920 14.560 35.840 14.840 ;
        RECT 0.000 14.280 4.200 14.560 ;
      LAYER met2 ;
        RECT 4.200 14.280 5.320 14.560 ;
      LAYER met2 ;
        RECT 5.320 14.280 5.880 14.560 ;
      LAYER met2 ;
        RECT 5.880 14.280 8.120 14.560 ;
      LAYER met2 ;
        RECT 8.120 14.280 9.240 14.560 ;
      LAYER met2 ;
        RECT 9.240 14.280 10.080 14.560 ;
      LAYER met2 ;
        RECT 10.080 14.280 24.360 14.560 ;
      LAYER met2 ;
        RECT 24.360 14.280 28.560 14.560 ;
      LAYER met2 ;
        RECT 28.560 14.280 30.520 14.560 ;
      LAYER met2 ;
        RECT 30.520 14.280 32.200 14.560 ;
      LAYER met2 ;
        RECT 32.200 14.280 35.840 14.560 ;
        RECT 0.000 13.720 3.920 14.280 ;
      LAYER met2 ;
        RECT 3.920 14.000 5.320 14.280 ;
      LAYER met2 ;
        RECT 5.320 14.000 5.600 14.280 ;
      LAYER met2 ;
        RECT 5.600 14.000 8.400 14.280 ;
      LAYER met2 ;
        RECT 8.400 14.000 8.960 14.280 ;
      LAYER met2 ;
        RECT 8.960 14.000 10.080 14.280 ;
        RECT 3.920 13.720 5.040 14.000 ;
      LAYER met2 ;
        RECT 0.000 13.160 3.640 13.720 ;
      LAYER met2 ;
        RECT 3.640 13.440 5.040 13.720 ;
      LAYER met2 ;
        RECT 5.040 13.440 5.600 14.000 ;
      LAYER met2 ;
        RECT 5.600 13.720 7.000 14.000 ;
      LAYER met2 ;
        RECT 7.000 13.720 7.280 14.000 ;
      LAYER met2 ;
        RECT 5.600 13.440 6.720 13.720 ;
      LAYER met2 ;
        RECT 6.720 13.440 7.280 13.720 ;
      LAYER met2 ;
        RECT 7.280 13.440 10.080 14.000 ;
      LAYER met2 ;
        RECT 10.080 13.720 24.080 14.280 ;
      LAYER met2 ;
        RECT 24.080 14.000 28.280 14.280 ;
      LAYER met2 ;
        RECT 28.280 14.000 30.800 14.280 ;
      LAYER met2 ;
        RECT 30.800 14.000 32.480 14.280 ;
        RECT 24.080 13.720 25.480 14.000 ;
      LAYER met2 ;
        RECT 25.480 13.720 25.760 14.000 ;
      LAYER met2 ;
        RECT 25.760 13.720 28.000 14.000 ;
      LAYER met2 ;
        RECT 28.000 13.720 31.080 14.000 ;
      LAYER met2 ;
        RECT 31.080 13.720 32.480 14.000 ;
      LAYER met2 ;
        RECT 32.480 13.720 35.840 14.280 ;
        RECT 10.080 13.440 20.720 13.720 ;
      LAYER met2 ;
        RECT 20.720 13.440 21.560 13.720 ;
      LAYER met2 ;
        RECT 21.560 13.440 24.080 13.720 ;
      LAYER met2 ;
        RECT 24.080 13.440 25.200 13.720 ;
      LAYER met2 ;
        RECT 25.200 13.440 25.760 13.720 ;
      LAYER met2 ;
        RECT 25.760 13.440 27.440 13.720 ;
      LAYER met2 ;
        RECT 27.440 13.440 31.360 13.720 ;
      LAYER met2 ;
        RECT 31.360 13.440 32.760 13.720 ;
      LAYER met2 ;
        RECT 32.760 13.440 35.840 13.720 ;
      LAYER met2 ;
        RECT 3.640 13.160 4.760 13.440 ;
      LAYER met2 ;
        RECT 0.000 10.640 3.360 13.160 ;
      LAYER met2 ;
        RECT 3.360 12.880 4.760 13.160 ;
      LAYER met2 ;
        RECT 4.760 12.880 7.560 13.440 ;
      LAYER met2 ;
        RECT 7.560 13.160 9.800 13.440 ;
      LAYER met2 ;
        RECT 9.800 13.160 17.080 13.440 ;
      LAYER met2 ;
        RECT 17.080 13.160 17.920 13.440 ;
      LAYER met2 ;
        RECT 17.920 13.160 20.160 13.440 ;
      LAYER met2 ;
        RECT 20.160 13.160 21.560 13.440 ;
        RECT 7.560 12.880 9.240 13.160 ;
      LAYER met2 ;
        RECT 9.240 12.880 16.800 13.160 ;
      LAYER met2 ;
        RECT 16.800 12.880 18.200 13.160 ;
      LAYER met2 ;
        RECT 18.200 12.880 19.880 13.160 ;
      LAYER met2 ;
        RECT 19.880 12.880 21.560 13.160 ;
      LAYER met2 ;
        RECT 21.560 12.880 25.760 13.440 ;
      LAYER met2 ;
        RECT 25.760 13.160 27.160 13.440 ;
      LAYER met2 ;
        RECT 27.160 13.160 31.640 13.440 ;
      LAYER met2 ;
        RECT 25.760 12.880 26.880 13.160 ;
      LAYER met2 ;
        RECT 26.880 12.880 31.640 13.160 ;
      LAYER met2 ;
        RECT 31.640 12.880 33.040 13.440 ;
      LAYER met2 ;
        RECT 33.040 12.880 35.840 13.440 ;
      LAYER met2 ;
        RECT 3.360 12.320 4.480 12.880 ;
      LAYER met2 ;
        RECT 4.480 12.600 16.520 12.880 ;
      LAYER met2 ;
        RECT 16.520 12.600 21.560 12.880 ;
      LAYER met2 ;
        RECT 21.560 12.600 31.920 12.880 ;
        RECT 4.480 12.320 14.000 12.600 ;
      LAYER met2 ;
        RECT 14.000 12.320 15.400 12.600 ;
      LAYER met2 ;
        RECT 15.400 12.320 15.960 12.600 ;
      LAYER met2 ;
        RECT 15.960 12.320 21.000 12.600 ;
      LAYER met2 ;
        RECT 21.000 12.320 31.920 12.600 ;
      LAYER met2 ;
        RECT 31.920 12.320 33.320 12.880 ;
        RECT 3.360 11.480 4.200 12.320 ;
      LAYER met2 ;
        RECT 4.200 11.760 14.000 12.320 ;
      LAYER met2 ;
        RECT 14.000 12.040 20.720 12.320 ;
      LAYER met2 ;
        RECT 20.720 12.040 31.360 12.320 ;
      LAYER met2 ;
        RECT 31.360 12.040 33.320 12.320 ;
      LAYER met2 ;
        RECT 33.320 12.040 35.840 12.880 ;
      LAYER met2 ;
        RECT 14.000 11.760 17.360 12.040 ;
      LAYER met2 ;
        RECT 17.360 11.760 18.200 12.040 ;
      LAYER met2 ;
        RECT 18.200 11.760 19.880 12.040 ;
      LAYER met2 ;
        RECT 19.880 11.760 26.880 12.040 ;
      LAYER met2 ;
        RECT 26.880 11.760 28.000 12.040 ;
      LAYER met2 ;
        RECT 28.000 11.760 30.800 12.040 ;
      LAYER met2 ;
        RECT 30.800 11.760 33.040 12.040 ;
      LAYER met2 ;
        RECT 33.040 11.760 35.840 12.040 ;
        RECT 4.200 11.480 14.560 11.760 ;
      LAYER met2 ;
        RECT 14.560 11.480 16.800 11.760 ;
      LAYER met2 ;
        RECT 16.800 11.480 26.600 11.760 ;
      LAYER met2 ;
        RECT 26.600 11.480 28.000 11.760 ;
      LAYER met2 ;
        RECT 28.000 11.480 29.120 11.760 ;
      LAYER met2 ;
        RECT 29.120 11.480 32.760 11.760 ;
      LAYER met2 ;
        RECT 32.760 11.480 35.840 11.760 ;
      LAYER met2 ;
        RECT 3.360 11.200 5.040 11.480 ;
      LAYER met2 ;
        RECT 5.040 11.200 6.440 11.480 ;
      LAYER met2 ;
        RECT 6.440 11.200 8.680 11.480 ;
      LAYER met2 ;
        RECT 8.680 11.200 26.320 11.480 ;
      LAYER met2 ;
        RECT 26.320 11.200 32.200 11.480 ;
      LAYER met2 ;
        RECT 32.200 11.200 35.840 11.480 ;
      LAYER met2 ;
        RECT 3.360 10.920 9.240 11.200 ;
      LAYER met2 ;
        RECT 9.240 10.920 25.760 11.200 ;
      LAYER met2 ;
        RECT 25.760 10.920 27.720 11.200 ;
      LAYER met2 ;
        RECT 27.720 10.920 28.000 11.200 ;
      LAYER met2 ;
        RECT 28.000 10.920 31.360 11.200 ;
      LAYER met2 ;
        RECT 31.360 10.920 35.840 11.200 ;
      LAYER met2 ;
        RECT 3.360 10.640 9.520 10.920 ;
      LAYER met2 ;
        RECT 9.520 10.640 25.200 10.920 ;
      LAYER met2 ;
        RECT 25.200 10.640 27.440 10.920 ;
      LAYER met2 ;
        RECT 27.440 10.640 28.000 10.920 ;
      LAYER met2 ;
        RECT 28.000 10.640 29.960 10.920 ;
      LAYER met2 ;
        RECT 29.960 10.640 35.840 10.920 ;
        RECT 0.000 10.360 4.200 10.640 ;
      LAYER met2 ;
        RECT 4.200 10.360 7.280 10.640 ;
      LAYER met2 ;
        RECT 7.280 10.360 7.840 10.640 ;
      LAYER met2 ;
        RECT 7.840 10.360 10.080 10.640 ;
      LAYER met2 ;
        RECT 10.080 10.360 24.640 10.640 ;
      LAYER met2 ;
        RECT 24.640 10.360 27.160 10.640 ;
      LAYER met2 ;
        RECT 27.160 10.360 35.840 10.640 ;
        RECT 0.000 10.080 8.400 10.360 ;
      LAYER met2 ;
        RECT 8.400 10.080 10.640 10.360 ;
      LAYER met2 ;
        RECT 10.640 10.080 23.800 10.360 ;
      LAYER met2 ;
        RECT 23.800 10.080 26.600 10.360 ;
      LAYER met2 ;
        RECT 26.600 10.080 35.840 10.360 ;
        RECT 0.000 9.800 8.680 10.080 ;
      LAYER met2 ;
        RECT 8.680 9.800 12.880 10.080 ;
      LAYER met2 ;
        RECT 12.880 9.800 22.960 10.080 ;
      LAYER met2 ;
        RECT 22.960 9.800 26.040 10.080 ;
      LAYER met2 ;
        RECT 26.040 9.800 35.840 10.080 ;
        RECT 0.000 9.520 9.240 9.800 ;
      LAYER met2 ;
        RECT 9.240 9.520 13.440 9.800 ;
      LAYER met2 ;
        RECT 13.440 9.520 22.960 9.800 ;
      LAYER met2 ;
        RECT 22.960 9.520 25.200 9.800 ;
      LAYER met2 ;
        RECT 25.200 9.520 35.840 9.800 ;
        RECT 0.000 9.240 9.800 9.520 ;
      LAYER met2 ;
        RECT 9.800 9.240 15.120 9.520 ;
      LAYER met2 ;
        RECT 15.120 9.240 22.960 9.520 ;
      LAYER met2 ;
        RECT 22.960 9.240 24.360 9.520 ;
      LAYER met2 ;
        RECT 24.360 9.240 35.840 9.520 ;
        RECT 0.000 8.680 10.360 9.240 ;
      LAYER met2 ;
        RECT 10.360 8.960 11.480 9.240 ;
      LAYER met2 ;
        RECT 11.480 8.960 12.040 9.240 ;
      LAYER met2 ;
        RECT 12.040 8.960 15.120 9.240 ;
      LAYER met2 ;
        RECT 15.120 8.960 35.840 9.240 ;
      LAYER met2 ;
        RECT 10.360 8.680 11.760 8.960 ;
      LAYER met2 ;
        RECT 11.760 8.680 12.880 8.960 ;
      LAYER met2 ;
        RECT 12.880 8.680 15.120 8.960 ;
      LAYER met2 ;
        RECT 15.120 8.680 24.080 8.960 ;
        RECT 0.000 8.120 10.640 8.680 ;
      LAYER met2 ;
        RECT 10.640 8.400 11.760 8.680 ;
      LAYER met2 ;
        RECT 11.760 8.400 24.080 8.680 ;
      LAYER met2 ;
        RECT 24.080 8.400 25.200 8.960 ;
      LAYER met2 ;
        RECT 25.200 8.400 35.840 8.960 ;
      LAYER met2 ;
        RECT 10.640 8.120 12.040 8.400 ;
      LAYER met2 ;
        RECT 12.040 8.120 24.080 8.400 ;
      LAYER met2 ;
        RECT 24.080 8.120 25.480 8.400 ;
      LAYER met2 ;
        RECT 25.480 8.120 35.840 8.400 ;
        RECT 0.000 7.560 10.920 8.120 ;
      LAYER met2 ;
        RECT 10.920 7.840 12.320 8.120 ;
      LAYER met2 ;
        RECT 12.320 7.840 24.360 8.120 ;
      LAYER met2 ;
        RECT 10.920 7.560 12.600 7.840 ;
      LAYER met2 ;
        RECT 12.600 7.560 24.360 7.840 ;
      LAYER met2 ;
        RECT 24.360 7.560 25.760 8.120 ;
      LAYER met2 ;
        RECT 0.000 7.280 11.200 7.560 ;
      LAYER met2 ;
        RECT 11.200 7.280 12.880 7.560 ;
      LAYER met2 ;
        RECT 12.880 7.280 24.640 7.560 ;
      LAYER met2 ;
        RECT 24.640 7.280 25.760 7.560 ;
      LAYER met2 ;
        RECT 25.760 7.280 35.840 8.120 ;
        RECT 0.000 7.000 11.480 7.280 ;
      LAYER met2 ;
        RECT 11.480 7.000 13.160 7.280 ;
      LAYER met2 ;
        RECT 0.000 6.720 11.760 7.000 ;
      LAYER met2 ;
        RECT 11.760 6.720 13.160 7.000 ;
      LAYER met2 ;
        RECT 13.160 6.720 24.920 7.280 ;
      LAYER met2 ;
        RECT 24.920 6.720 26.040 7.280 ;
      LAYER met2 ;
        RECT 26.040 6.720 35.840 7.280 ;
        RECT 0.000 6.440 12.040 6.720 ;
      LAYER met2 ;
        RECT 12.040 6.440 13.160 6.720 ;
      LAYER met2 ;
        RECT 0.000 5.880 11.760 6.440 ;
      LAYER met2 ;
        RECT 11.760 5.880 13.160 6.440 ;
      LAYER met2 ;
        RECT 13.160 5.880 25.200 6.720 ;
      LAYER met2 ;
        RECT 25.200 5.880 26.320 6.720 ;
      LAYER met2 ;
        RECT 0.000 5.600 11.480 5.880 ;
      LAYER met2 ;
        RECT 11.480 5.600 12.880 5.880 ;
      LAYER met2 ;
        RECT 12.880 5.600 25.480 5.880 ;
      LAYER met2 ;
        RECT 25.480 5.600 26.320 5.880 ;
      LAYER met2 ;
        RECT 26.320 5.600 35.840 6.720 ;
        RECT 0.000 5.320 11.200 5.600 ;
      LAYER met2 ;
        RECT 11.200 5.320 12.600 5.600 ;
      LAYER met2 ;
        RECT 12.600 5.320 25.480 5.600 ;
        RECT 0.000 5.040 10.920 5.320 ;
      LAYER met2 ;
        RECT 10.920 5.040 12.320 5.320 ;
      LAYER met2 ;
        RECT 0.000 3.920 10.640 5.040 ;
      LAYER met2 ;
        RECT 10.640 4.760 12.320 5.040 ;
      LAYER met2 ;
        RECT 12.320 4.760 25.480 5.320 ;
      LAYER met2 ;
        RECT 25.480 4.760 26.600 5.600 ;
      LAYER met2 ;
        RECT 26.600 4.760 35.840 5.600 ;
      LAYER met2 ;
        RECT 10.640 4.480 13.720 4.760 ;
      LAYER met2 ;
        RECT 13.720 4.480 25.760 4.760 ;
      LAYER met2 ;
        RECT 10.640 3.920 14.000 4.480 ;
      LAYER met2 ;
        RECT 14.000 3.920 25.760 4.480 ;
      LAYER met2 ;
        RECT 25.760 3.920 26.880 4.760 ;
      LAYER met2 ;
        RECT 0.000 3.080 12.600 3.920 ;
      LAYER met2 ;
        RECT 12.600 3.640 14.000 3.920 ;
      LAYER met2 ;
        RECT 14.000 3.640 26.040 3.920 ;
      LAYER met2 ;
        RECT 26.040 3.640 26.880 3.920 ;
      LAYER met2 ;
        RECT 26.880 3.640 35.840 4.760 ;
      LAYER met2 ;
        RECT 12.600 3.080 13.720 3.640 ;
      LAYER met2 ;
        RECT 13.720 3.080 26.040 3.640 ;
      LAYER met2 ;
        RECT 26.040 3.080 27.160 3.640 ;
      LAYER met2 ;
        RECT 0.000 2.240 12.320 3.080 ;
      LAYER met2 ;
        RECT 12.320 2.520 13.440 3.080 ;
      LAYER met2 ;
        RECT 13.440 2.520 26.320 3.080 ;
      LAYER met2 ;
        RECT 26.320 2.520 27.160 3.080 ;
      LAYER met2 ;
        RECT 27.160 2.520 35.840 3.640 ;
      LAYER met2 ;
        RECT 12.320 2.240 13.160 2.520 ;
      LAYER met2 ;
        RECT 0.000 0.280 12.040 2.240 ;
      LAYER met2 ;
        RECT 12.040 1.680 13.160 2.240 ;
      LAYER met2 ;
        RECT 13.160 1.680 26.320 2.520 ;
      LAYER met2 ;
        RECT 26.320 1.680 27.440 2.520 ;
        RECT 12.040 0.280 12.880 1.680 ;
      LAYER met2 ;
        RECT 12.880 0.280 26.600 1.680 ;
      LAYER met2 ;
        RECT 26.600 0.280 27.440 1.680 ;
      LAYER met2 ;
        RECT 27.440 0.280 35.840 2.520 ;
        RECT 0.000 0.000 35.840 0.280 ;
      LAYER met3 ;
        RECT 0.000 0.000 35.840 35.840 ;
      LAYER met4 ;
        RECT 0.000 0.000 35.840 35.840 ;
      LAYER met5 ;
        RECT 0.000 0.000 35.840 35.840 ;
  END
END my_logo
END LIBRARY

